
* Circuit Extracted by Tanner Research's L-Edit Version 15.00 / Extract Version 15.00 ;CMOSNuit Extracted by Tanner Research's L-Edit Version 15.00 / Extract Version 15.00 
* TDB File:  C:\Documents and Settings\Owner\Desktop\final\Layout_without_pads.tdb
* Cell:  Cell0	Version 1.87
* Extract Definition File:  mhp_n05.ext
* Extract Date and Time:  02/11/2022 - 01:15

* Tech: AMI_C5N
* LOT: T22Y_TT (typical)                  WAF: 3104
* Temperature_parameters=Optimized 
.MODEL CMOSN NMOS (                                LEVEL   = 7
+VERSION = 3.1            TNOM    = 27             TOX     = 1.39E-8
+XJ      = 1.5E-7         NCH     = 1.7E17         VTH0    = 0.6696061
+K1      = 0.8351612      K2      = -0.0839158     K3      = 23.1023856
+K3B     = -7.6841108     W0      = 1E-8           NLX     = 1E-9
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 2.9047241      DVT1    = 0.4302695      DVT2    = -0.134857
+U0      = 458.439679     UA      = 1E-13          UB      = 1.485499E-18
+UC      = 1.629939E-11   VSAT    = 1.643993E5     A0      = 0.6103537
+AGS     = 0.1194608      B0      = 2.674756E-6    B1      = 5E-6
+KETA    = -2.640681E-3   A1      = 8.219585E-5    A2      = 0.3564792
+RDSW    = 1.387108E3     PRWG    = 0.0299916      PRWB    = 0.0363981
+WR      = 1              WINT    = 2.472348E-7    LINT    = 3.597605E-8
+XL      = 0              XW      = 0              DWG     = -1.287163E-8
+DWB     = 5.306586E-8    VOFF    = 0              NFACTOR = 0.8365585
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 0.0246738      ETAB    = -1.406123E-3
+DSUB    = 0.2543458      PCLM    = 2.5945188      PDIBLC1 = -0.4282336
+PDIBLC2 = 2.311743E-3    PDIBLCB = -0.0272914     DROUT   = 0.7283566
+PSCBE1  = 5.598623E8     PSCBE2  = 5.461645E-5    PVAG    = 0
+DELTA   = 0.01           RSH     = 81.8           MOBMOD  = 1
+PRT     = 8.621          UTE     = -1             KT1     = -0.2501
+KT1L    = -2.58E-9       KT2     = 0              UA1     = 5.4E-10
+UB1     = -4.8E-19       UC1     = -7.5E-11       AT      = 1E5
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 2E-10          CGSO    = 2E-10          CGBO    = 1E-9
+CJ      = 4.197772E-4    PB      = 0.99           MJ      = 0.4515044
+CJSW    = 3.242724E-10   PBSW    = 0.1            MJSW    = 0.1153991
+CJSWG   = 1.64E-10       PBSWG   = 0.1            MJSWG   = 0.1153991
+CF      = 0              PVTH0   = 0.0585501      PRDSW   = 133.285505
+PK2     = -0.0299638     WKETA   = -0.0248758     LKETA   = 1.173187E-3
+AF      = 1              KF      = 0)
*
.MODEL CMOSP PMOS (                                LEVEL   = 7
+VERSION = 3.1            TNOM    = 27             TOX     = 1.39E-8
+XJ      = 1.5E-7         NCH     = 1.7E17         VTH0    = -0.9214347
+K1      = 0.5553722      K2      = 8.763328E-3    K3      = 6.3063558
+K3B     = -0.6487362     W0      = 1.280703E-8    NLX     = 2.593997E-8
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 2.5131165      DVT1    = 0.5480536      DVT2    = -0.1186489
+U0      = 212.0166131    UA      = 2.807115E-9    UB      = 1E-21
+UC      = -5.82128E-11   VSAT    = 1.713601E5     A0      = 0.8430019
+AGS     = 0.1328608      B0      = 7.117912E-7    B1      = 5E-6
+KETA    = -3.674859E-3   A1      = 4.77502E-5     A2      = 0.3
+RDSW    = 2.837206E3     PRWG    = -0.0363908     PRWB    = -1.016722E-5
+WR      = 1              WINT    = 2.838038E-7    LINT    = 5.528807E-8
+XL      = 0              XW      = 0              DWG     = -1.606385E-8
+DWB     = 2.266386E-8    VOFF    = -0.0558512     NFACTOR = 0.9342488
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 0.3251882      ETAB    = -0.0580325
+DSUB    = 1              PCLM    = 2.2409567      PDIBLC1 = 0.0411445
+PDIBLC2 = 3.355575E-3    PDIBLCB = -0.0551797     DROUT   = 0.2036901
+PSCBE1  = 6.44809E9      PSCBE2  = 6.300848E-10   PVAG    = 0
+DELTA   = 0.01           RSH     = 101.6          MOBMOD  = 1
+PRT     = 59.494         UTE     = -1             KT1     = -0.2942
+KT1L    = 1.68E-9        KT2     = 0              UA1     = 4.5E-9
+UB1     = -6.3E-18       UC1     = -1E-10         AT      = 1E3
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 2.9E-10        CGSO    = 2.9E-10        CGBO    = 1E-9
+CJ      = 7.235528E-4    PB      = 0.9527355      MJ      = 0.4955293
+CJSW    = 2.692786E-10   PBSW    = 0.99           MJSW    = 0.2958392
+CJSWG   = 6.4E-11        PBSWG   = 0.99           MJSWG   = 0.2958392
+CF      = 0              PVTH0   = 5.98016E-3     PRDSW   = 14.8598424
+PK2     = 3.73981E-3     WKETA   = 5.292165E-3    LKETA   = -4.205905E-3 
+AF      = 1              KF      = 0)
*

* Warning:  Layers with Unassigned FRINGE Capacitance.
*   <Pad Comment>

* NODE NAME ALIASES
*       10 = UAC34/U222/B (79.5 , 1259.5)
*       10 = UAC111/U223/vout (-1480 , 1258.5)
*       10 = UAC111/An (-1481 , 1302.5)
*       10 = UAC34/U206/A (136.5 , 1264.5)
*       10 = UAC34/A6 (138 , 1294)
*       11 = UAC34/U229/Vin (111 , 1217)
*       11 = UAC34/U220/OUT (109.5 , 1248)
*       12 = UAC111/U228/vout (-1388 , 1258.5)
*       12 = UAC111/D (-1351.5 , 1254)
*       12 = UAC111/Dn (-1389.5 , 1300.5)
*       12 = UAC31/D (-1205 , 1256)
*       12 = UAC31/U219/B (-1140.5 , 1259.5)
*       12 = UAC31/D6 (-1141 , 1286.5)
*       12 = UAC31/U220/B (-969 , 1259.5)
*       12 = UAC32/D (-841.5 , 1256)
*       12 = UAC32/U219/B (-777 , 1259.5)
*       12 = UAC32/D6 (-777.5 , 1286.5)
*       12 = UAC32/U220/B (-605.5 , 1259.5)
*       12 = UAC33/D (-477 , 1256)
*       12 = UAC33/U219/B (-412.5 , 1259.5)
*       12 = UAC33/D6 (-413 , 1286.5)
*       12 = UAC33/U220/B (-241 , 1259.5)
*       12 = UAC34/D (-113.5 , 1256)
*       12 = UAC34/U219/B (-49 , 1259.5)
*       12 = UAC34/D6 (-49.5 , 1286.5)
*       12 = UAC34/U220/B (122.5 , 1259.5)
*       19 = UAC34/U219/OUT (-62 , 1248)
*       19 = UAC34/U262/vin (-12 , 1260)
*       20 = UAC34/U262/vout (-26.5 , 1261.5)
*       20 = UAC34/U222/A (6 , 1264.5)
*       27 = UAC33/U206/Vout (-191.5 , 1271.5)
*       27 = UAC33/U236/A (-168.5 , 1215.5)
*       27 = UAC33/U235/B (-186.5 , 1215.5)
*       35 = UAC33/U218/B (-277.5 , 1215.5)
*       35 = UAC33/U229/Vout (-238.5 , 1217)
*       39 = UAC33/U219/OUT (-425.5 , 1248)
*       39 = UAC33/U262/vin (-375.5 , 1260)
*       40 = UAC33/U222/A (-357.5 , 1264.5)
*       40 = UAC33/U262/vout (-390 , 1261.5)
*       56 = UAC32/U262/vout (-754.5 , 1261.5)
*       56 = UAC32/U222/A (-722 , 1264.5)
*       58 = UAC32/U219/OUT (-790 , 1248)
*       58 = UAC32/U262/vin (-740 , 1260)
*       65 = UAC111/U220/B (-1387 , 1169)
*       65 = UAC111/U230/vout (-1367 , 1213)
*       65 = UAC111/Fn (-1351 , 1237)
*       65 = UAC31/F (-1205 , 1268)
*       65 = UAC32/F (-841.5 , 1268)
*       65 = UAC31/U206/B (-881.5 , 1259.5)
*       65 = UAC31/F6 (-877.5 , 1288)
*       65 = UAC32/U206/B (-518 , 1259.5)
*       65 = UAC32/F6 (-514 , 1288)
*       65 = UAC33/F (-477 , 1268)
*       65 = UAC34/F (-113.5 , 1268)
*       65 = UAC33/U206/B (-153.5 , 1259.5)
*       65 = UAC33/F6 (-149.5 , 1288)
*       65 = UAC34/U206/B (210 , 1259.5)
*       65 = UAC34/F6 (214 , 1288)
*       71 = UAC31/U238/B (-1141 , 1215.5)
*       71 = UAC31/U220/A (-995.5 , 1259.5)
*       71 = UAC31/C6 (-995.5 , 1291.5)
*       71 = UAC32/U254/Vout (-673 , 1173)
*       71 = UAC32/P (-672 , 1146)
*       71 = UAC31/U236/B (-870 , 1215.5)
*       71 = UAC31/C (-829.5 , 1242.5)
*       77 = UAC31/U219/OUT (-1153.5 , 1248)
*       77 = UAC31/U262/vin (-1103.5 , 1260)
*       78 = UAC31/U262/vout (-1118 , 1261.5)
*       78 = UAC31/U222/A (-1085.5 , 1264.5)
*       80 = UAC111/U228/vin (-1416.5 , 1259.5)
*       80 = UAC111/U227/O/P (-1432 , 1267.5)
*       82 = UAC111/U223/vin (-1508.5 , 1259.5)
*       82 = UAC111/U222/OUT (-1539 , 1248)
*       84 = UAC34/U246/Vin (203 , 1173)
*       84 = UAC34/U236/OUT (208.5 , 1204)
*       85 = UAC34/U253/C (125 , 1161.5)
*       85 = UAC34/U247/Vout (169 , 1173)
*       86 = UAC34/U247/Vin (155 , 1173)
*       86 = UAC34/U235/OUT (164 , 1204)
*       87 = UAC34/U236/A (195 , 1215.5)
*       87 = UAC34/U235/B (177 , 1215.5)
*       87 = UAC34/U206/Vout (172 , 1271.5)
*       88 = UAC34/U236/VDD (200.5 , 1237)
*       88 = UAC34/U235/VDD (156 , 1237)
*       88 = UAC34/U229/Vdd (119 , 1237.5)
*       88 = UAC34/U245/Vdd (-15 , 1237.5)
*       88 = UAC34/U238/VDD (-70.5 , 1237)
*       88 = UAC34/U218/VDD (9 , 1234.5)
*       88 = UAC34/U220/VDD (101.5 , 1281)
*       88 = UAC33/U238/VDD (-434 , 1237)
*       88 = UAC33/U245/Vdd (-378.5 , 1237.5)
*       88 = UAC33/U218/VDD (-354.5 , 1234.5)
*       88 = UAC33/U235/VDD (-207.5 , 1237)
*       88 = UAC33/U229/Vdd (-244.5 , 1237.5)
*       88 = UAC33/U222/VDD (-361 , 1278.5)
*       88 = UAC32/U238/VDD (-798.5 , 1237)
*       88 = UAC32/U245/Vdd (-743 , 1237.5)
*       88 = UAC32/U218/VDD (-719 , 1234.5)
*       88 = UAC32/U229/Vdd (-609 , 1237.5)
*       88 = UAC32/U236/VDD (-527.5 , 1237)
*       88 = UAC32/U235/VDD (-572 , 1237)
*       88 = UAC32/U206/VDD (-591.002 , 1278.5)
*       88 = UAC31/U245/Vdd (-1106.5 , 1237.5)
*       88 = UAC31/U238/VDD (-1162 , 1237)
*       88 = UAC31/U218/VDD (-1082.5 , 1234.5)
*       88 = UAC31/U235/VDD (-935.5 , 1237)
*       88 = UAC31/U229/Vdd (-972.5 , 1237.5)
*       88 = UAC31/U206/VDD (-958.5 , 1278.5)
*       88 = UAC31/U220/VDD (-990 , 1281)
*       88 = UAC111/U225/VDD (-1518 , 1235.5)
*       88 = UAC111/U224/Vdd (-1554 , 1236.5)
*       88 = UAC111/U223/Vdd (-1499 , 1282)
*       88 = UAC111/U222/VDD (-1547 , 1281)
*       88 = UAC111/U231/VDD (-1539 , 1190.5)
*       88 = UAC111/U220/VDD (-1464 , 1188)
*       88 = UAC111/U232/Vdd (-1491 , 1191.5)
*       88 = UAC111/U229/VDD (-1434 , 1235.5)
*       88 = UAC111/U226/Vdd (-1470 , 1236.5)
*       88 = UAC111/Fn (-1591 , 1225.5)
*       88 = UAC111/U229/B (-1413 , 1214)
*       88 = UAC111/U228/Vdd (-1407 , 1282)
*       88 = UAC111/U227/VDD (-1425.5 , 1279.5)
*       88 = UAC111/F (-1409.5 , 1299.5)
*       88 = UAC111/U230/Vdd (-1386 , 1236.5)
*       88 = UAC31/U262/VDD (-1125 , 1282)
*       88 = UAC31/U219/VDD (-1161.5 , 1281)
*       88 = UAC31/U222/VDD (-1089 , 1278.5)
*       88 = UAC32/U219/VDD (-798 , 1281)
*       88 = UAC31/U236/VDD (-891 , 1237)
*       88 = UAC31/U254/Vdd (-1042.5 , 1193.5)
*       88 = UAC31/U253/VDD (-956.5 , 1191.5)
*       88 = UAC31/U247/Vdd (-928.5 , 1193.5)
*       88 = UAC31/U246/Vdd (-880.5 , 1193.5)
*       88 = UAC32/U262/VDD (-761.5 , 1282)
*       88 = UAC32/U222/VDD (-725.5 , 1278.5)
*       88 = UAC32/U220/VDD (-626.5 , 1281)
*       88 = UAC32/U254/Vdd (-679 , 1193.5)
*       88 = UAC32/U253/VDD (-593 , 1191.5)
*       88 = UAC32/U247/Vdd (-565 , 1193.5)
*       88 = UAC32/U246/Vdd (-517 , 1193.5)
*       88 = UAC33/U262/VDD (-397 , 1282)
*       88 = UAC33/U219/VDD (-433.5 , 1281)
*       88 = UAC33/U206/VDD (-230.5 , 1278.5)
*       88 = UAC33/U220/VDD (-262 , 1281)
*       88 = UAC33/U236/VDD (-163 , 1237)
*       88 = UAC33/U254/Vdd (-314.5 , 1193.5)
*       88 = UAC33/U253/VDD (-228.5 , 1191.5)
*       88 = UAC33/U247/Vdd (-200.5 , 1193.5)
*       88 = UAC33/U246/Vdd (-152.5 , 1193.5)
*       88 = UAC34/U262/VDD (-33.5 , 1282)
*       88 = UAC34/U222/VDD (2.5 , 1278.5)
*       88 = UAC34/U219/VDD (-70 , 1281)
*       88 = UAC34/U206/VDD (133 , 1278.5)
*       88 = UAC34/U254/Vdd (49 , 1193.5)
*       88 = UAC34/U253/VDD (135 , 1191.5)
*       88 = UAC34/U247/Vdd (163 , 1193.5)
*       88 = UAC38/U245/Vdd (-15.5 , 1075)
*       88 = UAC38/U238/VDD (-71 , 1074.5)
*       88 = UAC38/U218/VDD (8.5 , 1072)
*       88 = UAC38/U236/VDD (200 , 1074.5)
*       88 = UAC38/U235/VDD (155.5 , 1074.5)
*       88 = UAC38/U229/Vdd (118.5 , 1075)
*       88 = UAC38/U220/VDD (101 , 1118.5)
*       88 = UAC37/U238/VDD (-434.5 , 1074.5)
*       88 = UAC37/U245/Vdd (-379 , 1075)
*       88 = UAC37/U218/VDD (-355 , 1072)
*       88 = UAC37/U235/VDD (-208 , 1074.5)
*       88 = UAC37/U229/Vdd (-245 , 1075)
*       88 = UAC37/U222/VDD (-361.5 , 1116)
*       88 = UAC36/U254/Vdd (-679.5 , 1031)
*       88 = UAC36/U253/VDD (-593.5 , 1029)
*       88 = UAC36/U247/Vdd (-565.5 , 1031)
*       88 = UAC36/U246/Vdd (-517.5 , 1031)
*       88 = UAC36/U238/VDD (-799 , 1074.5)
*       88 = UAC36/U245/Vdd (-743.5 , 1075)
*       88 = UAC36/U218/VDD (-719.5 , 1072)
*       88 = UAC36/U229/Vdd (-609.5 , 1075)
*       88 = UAC36/U236/VDD (-528 , 1074.5)
*       88 = UAC36/U235/VDD (-572.5 , 1074.5)
*       88 = UAC36/U206/VDD (-591.002 , 1116)
*       88 = UAC36/U219/VDD (-798.5 , 1118.5)
*       88 = UAC35/U246/Vdd (-881 , 1031)
*       88 = UAC35/U236/VDD (-891.5 , 1074.5)
*       88 = UAC35/U235/VDD (-936 , 1074.5)
*       88 = UAC35/U229/Vdd (-973 , 1075)
*       88 = UAC35/U245/Vdd (-1107 , 1075)
*       88 = UAC35/U238/VDD (-1162.5 , 1074.5)
*       88 = UAC35/U218/VDD (-1083 , 1072)
*       88 = UAC35/U206/VDD (-959 , 1116)
*       88 = UAC35/U220/VDD (-990.5 , 1118.5)
*       88 = UAC78/U245/Vdd (-1471 , 1075)
*       88 = UAC78/U218/VDD (-1447 , 1072)
*       88 = UAC78/U238/VDD (-1526.5 , 1074.5)
*       88 = UAC78/U235/VDD (-1300 , 1074.5)
*       88 = UAC78/U229/Vdd (-1337 , 1075)
*       88 = UAC112/U231/VDD (-1904.5 , 1028)
*       88 = UAC112/U224/Vdd (-1919.5 , 1074)
*       88 = UAC112/U222/VDD (-1912.5 , 1118.5)
*       88 = UAC112/U220/VDD (-1829.5 , 1025.5)
*       88 = UAC112/U232/Vdd (-1856.5 , 1029)
*       88 = UAC112/U229/VDD (-1799.5 , 1073)
*       88 = UAC112/U226/Vdd (-1835.5 , 1074)
*       88 = UAC112/U225/VDD (-1883.5 , 1073)
*       88 = UAC112/U223/Vdd (-1864.5 , 1119.5)
*       88 = UAC112/U230/Vdd (-1751.5 , 1074)
*       88 = UAC112/U228/Vdd (-1772.5 , 1119.5)
*       88 = UAC112/U227/VDD (-1791 , 1117)
*       88 = UAC78/U219/VDD (-1526 , 1118.5)
*       88 = UAC78/U262/VDD (-1489.5 , 1119.5)
*       88 = UAC78/U222/VDD (-1453.5 , 1116)
*       88 = UAC78/U206/VDD (-1323 , 1116)
*       88 = UAC78/U220/VDD (-1354.5 , 1118.5)
*       88 = UAC78/U254/Vdd (-1407 , 1031)
*       88 = UAC78/U253/VDD (-1321 , 1029)
*       88 = UAC78/U247/Vdd (-1293 , 1031)
*       88 = UAC78/U246/Vdd (-1245 , 1031)
*       88 = UAC78/U236/VDD (-1255.5 , 1074.5)
*       88 = UAC35/U262/VDD (-1125.5 , 1119.5)
*       88 = UAC35/U219/VDD (-1162 , 1118.5)
*       88 = UAC35/U222/VDD (-1089.5 , 1116)
*       88 = UAC35/U254/Vdd (-1043 , 1031)
*       88 = UAC35/U253/VDD (-957 , 1029)
*       88 = UAC35/U247/Vdd (-929 , 1031)
*       88 = UAC36/U262/VDD (-762 , 1119.5)
*       88 = UAC36/U222/VDD (-726 , 1116)
*       88 = UAC36/U220/VDD (-627 , 1118.5)
*       88 = UAC37/U262/VDD (-397.5 , 1119.5)
*       88 = UAC37/U219/VDD (-434 , 1118.5)
*       88 = UAC37/U206/VDD (-231 , 1116)
*       88 = UAC37/U220/VDD (-262.5 , 1118.5)
*       88 = UAC37/U254/Vdd (-315 , 1031)
*       88 = UAC37/U253/VDD (-229 , 1029)
*       88 = UAC37/U247/Vdd (-201 , 1031)
*       88 = UAC37/U246/Vdd (-153 , 1031)
*       88 = UAC37/U236/VDD (-163.5 , 1074.5)
*       88 = UAC38/U262/VDD (-34 , 1119.5)
*       88 = UAC38/U222/VDD (2 , 1116)
*       88 = UAC38/U219/VDD (-70.5 , 1118.5)
*       88 = UAC38/U206/VDD (132.5 , 1116)
*       88 = UAC42/U220/VDD (100.5 , 956)
*       88 = UAC41/U222/VDD (-362 , 953.5)
*       88 = UAC40/U206/VDD (-591.002 , 953.5)
*       88 = UAC39/U206/VDD (-959.5 , 953.5)
*       88 = UAC39/U220/VDD (-991 , 956)
*       88 = UAC80/U220/VDD (-1718.5 , 956)
*       88 = UAC80/U262/VDD (-1853.5 , 957)
*       88 = UAC80/U222/VDD (-1817.5 , 953.5)
*       88 = UAC80/U219/VDD (-1890 , 956)
*       88 = UAC114/U223/Vdd (-2241.5 , 957)
*       88 = UAC114/U222/VDD (-2289.5 , 956)
*       88 = UAC114/U220/VDD (-2206.5 , 863)
*       88 = UAC114/U232/Vdd (-2233.5 , 866.5)
*       88 = UAC114/U231/VDD (-2281.5 , 865.5)
*       88 = UAC114/U224/Vdd (-2296.5 , 911.5)
*       88 = UAC114/U226/Vdd (-2212.5 , 911.5)
*       88 = UAC114/U225/VDD (-2260.5 , 910.5)
*       88 = UAC114/U230/Vdd (-2128.5 , 911.5)
*       88 = UAC114/U229/VDD (-2176.5 , 910.5)
*       88 = UAC114/U228/Vdd (-2149.5 , 957)
*       88 = UAC114/U227/VDD (-2168 , 954.5)
*       88 = UAC80/U206/VDD (-1687 , 953.5)
*       88 = UAC80/U254/Vdd (-1771 , 868.5)
*       88 = UAC80/U253/VDD (-1685 , 866.5)
*       88 = UAC80/U247/Vdd (-1657 , 868.5)
*       88 = UAC80/U246/Vdd (-1609 , 868.5)
*       88 = UAC80/U245/Vdd (-1835 , 912.5)
*       88 = UAC80/U238/VDD (-1890.5 , 912)
*       88 = UAC80/U218/VDD (-1811 , 909.5)
*       88 = UAC80/U229/Vdd (-1701 , 912.5)
*       88 = UAC80/U236/VDD (-1619.5 , 912)
*       88 = UAC80/U235/VDD (-1664 , 912)
*       88 = UAC79/U219/VDD (-1526.5 , 956)
*       88 = UAC79/U262/VDD (-1490 , 957)
*       88 = UAC79/U222/VDD (-1454 , 953.5)
*       88 = UAC79/U206/VDD (-1323.5 , 953.5)
*       88 = UAC79/U220/VDD (-1355 , 956)
*       88 = UAC79/U245/Vdd (-1471.5 , 912.5)
*       88 = UAC79/U218/VDD (-1447.5 , 909.5)
*       88 = UAC79/U238/VDD (-1527 , 912)
*       88 = UAC79/U235/VDD (-1300.5 , 912)
*       88 = UAC79/U229/Vdd (-1337.5 , 912.5)
*       88 = UAC79/U254/Vdd (-1407.5 , 868.5)
*       88 = UAC79/U253/VDD (-1321.5 , 866.5)
*       88 = UAC79/U247/Vdd (-1293.5 , 868.5)
*       88 = UAC79/U246/Vdd (-1245.5 , 868.5)
*       88 = UAC79/U236/VDD (-1256 , 912)
*       88 = UAC39/U262/VDD (-1126 , 957)
*       88 = UAC39/U219/VDD (-1162.5 , 956)
*       88 = UAC39/U222/VDD (-1090 , 953.5)
*       88 = UAC39/U246/Vdd (-881.5 , 868.5)
*       88 = UAC39/U254/Vdd (-1043.5 , 868.5)
*       88 = UAC39/U253/VDD (-957.5 , 866.5)
*       88 = UAC39/U247/Vdd (-929.5 , 868.5)
*       88 = UAC39/U245/Vdd (-1107.5 , 912.5)
*       88 = UAC39/U238/VDD (-1163 , 912)
*       88 = UAC39/U218/VDD (-1083.5 , 909.5)
*       88 = UAC39/U236/VDD (-892 , 912)
*       88 = UAC39/U235/VDD (-936.5 , 912)
*       88 = UAC39/U229/Vdd (-973.5 , 912.5)
*       88 = UAC40/U219/VDD (-799 , 956)
*       88 = UAC40/U262/VDD (-762.5 , 957)
*       88 = UAC40/U222/VDD (-726.5 , 953.5)
*       88 = UAC40/U220/VDD (-627.5 , 956)
*       88 = UAC40/U254/Vdd (-680 , 868.5)
*       88 = UAC40/U253/VDD (-594 , 866.5)
*       88 = UAC40/U238/VDD (-799.5 , 912)
*       88 = UAC40/U245/Vdd (-744 , 912.5)
*       88 = UAC40/U218/VDD (-720 , 909.5)
*       88 = UAC40/U229/Vdd (-610 , 912.5)
*       88 = UAC40/U247/Vdd (-566 , 868.5)
*       88 = UAC40/U246/Vdd (-518 , 868.5)
*       88 = UAC40/U236/VDD (-528.5 , 912)
*       88 = UAC40/U235/VDD (-573 , 912)
*       88 = UAC41/U262/VDD (-398 , 957)
*       88 = UAC41/U219/VDD (-434.5 , 956)
*       88 = UAC41/U206/VDD (-231.5 , 953.5)
*       88 = UAC41/U220/VDD (-263 , 956)
*       88 = UAC41/U238/VDD (-435 , 912)
*       88 = UAC41/U245/Vdd (-379.5 , 912.5)
*       88 = UAC41/U218/VDD (-355.5 , 909.5)
*       88 = UAC41/U235/VDD (-208.5 , 912)
*       88 = UAC41/U229/Vdd (-245.5 , 912.5)
*       88 = UAC41/U254/Vdd (-315.5 , 868.5)
*       88 = UAC41/U253/VDD (-229.5 , 866.5)
*       88 = UAC41/U247/Vdd (-201.5 , 868.5)
*       88 = UAC41/U246/Vdd (-153.5 , 868.5)
*       88 = UAC41/U236/VDD (-164 , 912)
*       88 = UAC42/U262/VDD (-34.5 , 957)
*       88 = UAC42/U222/VDD (1.5 , 953.5)
*       88 = UAC42/U219/VDD (-71 , 956)
*       88 = UAC42/U206/VDD (132 , 953.5)
*       88 = UAC42/U254/Vdd (48 , 868.5)
*       88 = UAC42/U253/VDD (134 , 866.5)
*       88 = UAC42/U247/Vdd (162 , 868.5)
*       88 = UAC42/U245/Vdd (-16 , 912.5)
*       88 = UAC42/U238/VDD (-71.5 , 912)
*       88 = UAC42/U218/VDD (8 , 909.5)
*       88 = UAC42/U236/VDD (199.5 , 912)
*       88 = UAC42/U235/VDD (155 , 912)
*       88 = UAC42/U229/Vdd (118 , 912.5)
*       88 = UAC54/U236/VDD (199 , 750.5)
*       88 = UAC54/U235/VDD (154.5 , 750.5)
*       88 = UAC54/U229/Vdd (117.5 , 751)
*       88 = UAC54/U245/Vdd (-16.5 , 751)
*       88 = UAC54/U238/VDD (-72 , 750.5)
*       88 = UAC54/U218/VDD (7.5 , 748)
*       88 = UAC54/U220/VDD (100 , 794.5)
*       88 = UAC53/U238/VDD (-435.5 , 750.5)
*       88 = UAC53/U245/Vdd (-380 , 751)
*       88 = UAC53/U218/VDD (-356 , 748)
*       88 = UAC53/U235/VDD (-209 , 750.5)
*       88 = UAC53/U229/Vdd (-246 , 751)
*       88 = UAC53/U222/VDD (-362.5 , 792)
*       88 = UAC52/U206/VDD (-591.002 , 792)
*       88 = UAC52/U236/VDD (-529 , 750.5)
*       88 = UAC52/U235/VDD (-573.5 , 750.5)
*       88 = UAC52/U238/VDD (-800 , 750.5)
*       88 = UAC52/U245/Vdd (-744.5 , 751)
*       88 = UAC52/U218/VDD (-720.5 , 748)
*       88 = UAC52/U229/Vdd (-610.5 , 751)
*       88 = UAC51/U245/Vdd (-1108 , 751)
*       88 = UAC51/U238/VDD (-1163.5 , 750.5)
*       88 = UAC51/U218/VDD (-1084 , 748)
*       88 = UAC51/U236/VDD (-892.5 , 750.5)
*       88 = UAC51/U235/VDD (-937 , 750.5)
*       88 = UAC51/U229/Vdd (-974 , 751)
*       88 = UAC51/U206/VDD (-960 , 792)
*       88 = UAC81/U238/VDD (-1535 , 750.5)
*       88 = UAC81/U245/Vdd (-1479.5 , 751)
*       88 = UAC81/U218/VDD (-1455.5 , 748)
*       88 = UAC81/U235/VDD (-1308.5 , 750.5)
*       88 = UAC81/U229/Vdd (-1345.5 , 751)
*       88 = UAC81/U222/VDD (-1462 , 792)
*       88 = UAC82/U236/VDD (-1632.5 , 750.5)
*       88 = UAC82/U235/VDD (-1677 , 750.5)
*       88 = UAC82/U238/VDD (-1903.5 , 750.5)
*       88 = UAC82/U245/Vdd (-1848 , 751)
*       88 = UAC82/U218/VDD (-1824 , 748)
*       88 = UAC82/U229/Vdd (-1714 , 751)
*       88 = UAC84/U245/Vdd (-2211.5 , 751)
*       88 = UAC84/U238/VDD (-2267 , 750.5)
*       88 = UAC84/U218/VDD (-2187.5 , 748)
*       88 = UAC84/U236/VDD (-1996 , 750.5)
*       88 = UAC84/U235/VDD (-2040.5 , 750.5)
*       88 = UAC84/U229/Vdd (-2077.5 , 751)
*       88 = UAC116/U230/Vdd (-2499.5 , 750)
*       88 = UAC116/U229/VDD (-2547.5 , 749)
*       88 = UAC116/U226/Vdd (-2583.5 , 750)
*       88 = UAC116/U232/Vdd (-2604.5 , 705)
*       88 = UAC116/U231/VDD (-2652.5 , 704)
*       88 = UAC116/U220/VDD (-2577.5 , 701.5)
*       88 = UAC116/U225/VDD (-2631.5 , 749)
*       88 = UAC116/U224/Vdd (-2667.5 , 750)
*       88 = UAC116/U223/Vdd (-2612.5 , 795.5)
*       88 = UAC116/U222/VDD (-2660.5 , 794.5)
*       88 = UAC116/U228/Vdd (-2520.5 , 795.5)
*       88 = UAC116/U227/VDD (-2539 , 793)
*       88 = UAC84/U262/VDD (-2230 , 795.5)
*       88 = UAC84/U222/VDD (-2194 , 792)
*       88 = UAC84/U219/VDD (-2266.5 , 794.5)
*       88 = UAC84/U220/VDD (-2095 , 794.5)
*       88 = UAC84/U206/VDD (-2063.5 , 792)
*       88 = UAC84/U254/Vdd (-2147.5 , 707)
*       88 = UAC84/U253/VDD (-2061.5 , 705)
*       88 = UAC84/U247/Vdd (-2033.5 , 707)
*       88 = UAC84/U246/Vdd (-1985.5 , 707)
*       88 = UAC82/U219/VDD (-1903 , 794.5)
*       88 = UAC82/U262/VDD (-1866.5 , 795.5)
*       88 = UAC82/U222/VDD (-1830.5 , 792)
*       88 = UAC82/U206/VDD (-1700 , 792)
*       88 = UAC82/U220/VDD (-1731.5 , 794.5)
*       88 = UAC82/U254/Vdd (-1784 , 707)
*       88 = UAC82/U253/VDD (-1698 , 705)
*       88 = UAC82/U247/Vdd (-1670 , 707)
*       88 = UAC82/U246/Vdd (-1622 , 707)
*       88 = UAC81/U262/VDD (-1498 , 795.5)
*       88 = UAC81/U219/VDD (-1534.5 , 794.5)
*       88 = UAC81/U206/VDD (-1331.5 , 792)
*       88 = UAC81/U220/VDD (-1363 , 794.5)
*       88 = UAC81/U254/Vdd (-1415.5 , 707)
*       88 = UAC81/U253/VDD (-1329.5 , 705)
*       88 = UAC81/U247/Vdd (-1301.5 , 707)
*       88 = UAC81/U246/Vdd (-1253.5 , 707)
*       88 = UAC81/U236/VDD (-1264 , 750.5)
*       88 = UAC51/U262/VDD (-1126.5 , 795.5)
*       88 = UAC51/U219/VDD (-1163 , 794.5)
*       88 = UAC51/U222/VDD (-1090.5 , 792)
*       88 = UAC51/U220/VDD (-991.5 , 794.5)
*       88 = UAC51/U254/Vdd (-1044 , 707)
*       88 = UAC51/U253/VDD (-958 , 705)
*       88 = UAC51/U247/Vdd (-930 , 707)
*       88 = UAC51/U246/Vdd (-882 , 707)
*       88 = UAC52/U219/VDD (-799.5 , 794.5)
*       88 = UAC52/U262/VDD (-763 , 795.5)
*       88 = UAC52/U222/VDD (-727 , 792)
*       88 = UAC52/U220/VDD (-628 , 794.5)
*       88 = UAC52/U254/Vdd (-680.5 , 707)
*       88 = UAC52/U253/VDD (-594.5 , 705)
*       88 = UAC52/U247/Vdd (-566.5 , 707)
*       88 = UAC52/U246/Vdd (-518.5 , 707)
*       88 = UAC53/U262/VDD (-398.5 , 795.5)
*       88 = UAC53/U219/VDD (-435 , 794.5)
*       88 = UAC53/U206/VDD (-232 , 792)
*       88 = UAC53/U220/VDD (-263.5 , 794.5)
*       88 = UAC53/U254/Vdd (-316 , 707)
*       88 = UAC53/U253/VDD (-230 , 705)
*       88 = UAC53/U247/Vdd (-202 , 707)
*       88 = UAC53/U246/Vdd (-154 , 707)
*       88 = UAC53/U236/VDD (-164.5 , 750.5)
*       88 = UAC54/U262/VDD (-35 , 795.5)
*       88 = UAC54/U222/VDD (1 , 792)
*       88 = UAC54/U219/VDD (-71.5 , 794.5)
*       88 = UAC54/U206/VDD (131.5 , 792)
*       88 = UAC87/U254/Vdd (-1784 , 544.5)
*       88 = UAC87/U253/VDD (-1698 , 542.5)
*       88 = UAC87/U238/VDD (-1903.5 , 588)
*       88 = UAC87/U245/Vdd (-1848 , 588.5)
*       88 = UAC87/U218/VDD (-1824 , 585.5)
*       88 = UAC87/U229/Vdd (-1714 , 588.5)
*       88 = UAC87/U247/Vdd (-1670 , 544.5)
*       88 = UAC87/U246/Vdd (-1622 , 544.5)
*       88 = UAC87/U236/VDD (-1632.5 , 588)
*       88 = UAC87/U235/VDD (-1677 , 588)
*       88 = UAC118/U231/VDD (-3018.5 , 541.5)
*       88 = UAC118/U225/VDD (-2997.5 , 586.5)
*       88 = UAC118/U224/Vdd (-3033.5 , 587.5)
*       88 = UAC118/U220/VDD (-2943.5 , 539)
*       88 = UAC118/U232/Vdd (-2970.5 , 542.5)
*       88 = UAC118/U229/VDD (-2913.5 , 586.5)
*       88 = UAC118/U226/Vdd (-2949.5 , 587.5)
*       88 = UAC118/U230/Vdd (-2865.5 , 587.5)
*       88 = UAC118/U222/VDD (-3026.5 , 632)
*       88 = UAC118/U227/VDD (-2905 , 630.5)
*       88 = UAC118/U223/Vdd (-2978.5 , 633)
*       88 = UAC118/U228/Vdd (-2886.5 , 633)
*       88 = UAC90/U262/VDD (-2601 , 633)
*       88 = UAC90/U219/VDD (-2637.5 , 632)
*       88 = UAC90/U222/VDD (-2565 , 629.5)
*       88 = UAC90/U206/VDD (-2434.5 , 629.5)
*       88 = UAC90/U220/VDD (-2466 , 632)
*       88 = UAC90/U245/Vdd (-2582.5 , 588.5)
*       88 = UAC90/U218/VDD (-2558.5 , 585.5)
*       88 = UAC90/U238/VDD (-2638 , 588)
*       88 = UAC90/U235/VDD (-2411.5 , 588)
*       88 = UAC90/U229/Vdd (-2448.5 , 588.5)
*       88 = UAC90/U254/Vdd (-2518.5 , 544.5)
*       88 = UAC90/U253/VDD (-2432.5 , 542.5)
*       88 = UAC90/U247/Vdd (-2404.5 , 544.5)
*       88 = UAC90/U246/Vdd (-2356.5 , 544.5)
*       88 = UAC90/U236/VDD (-2367 , 588)
*       88 = UAC88/U262/VDD (-2230.5 , 633)
*       88 = UAC88/U222/VDD (-2194.5 , 629.5)
*       88 = UAC88/U219/VDD (-2267 , 632)
*       88 = UAC88/U220/VDD (-2095.5 , 632)
*       88 = UAC88/U206/VDD (-2064 , 629.5)
*       88 = UAC88/U254/Vdd (-2148 , 544.5)
*       88 = UAC88/U253/VDD (-2062 , 542.5)
*       88 = UAC88/U247/Vdd (-2034 , 544.5)
*       88 = UAC88/U245/Vdd (-2212 , 588.5)
*       88 = UAC88/U238/VDD (-2267.5 , 588)
*       88 = UAC88/U218/VDD (-2188 , 585.5)
*       88 = UAC88/U236/VDD (-1996.5 , 588)
*       88 = UAC88/U235/VDD (-2041 , 588)
*       88 = UAC88/U229/Vdd (-2078 , 588.5)
*       88 = UAC88/U246/Vdd (-1986 , 544.5)
*       88 = UAC87/U219/VDD (-1903 , 632)
*       88 = UAC87/U262/VDD (-1866.5 , 633)
*       88 = UAC87/U222/VDD (-1830.5 , 629.5)
*       88 = UAC87/U206/VDD (-1700 , 629.5)
*       88 = UAC87/U220/VDD (-1731.5 , 632)
*       88 = UAC85/U262/VDD (-1498.5 , 633)
*       88 = UAC85/U219/VDD (-1535 , 632)
*       88 = UAC85/U222/VDD (-1462.5 , 629.5)
*       88 = UAC85/U206/VDD (-1332 , 629.5)
*       88 = UAC85/U220/VDD (-1363.5 , 632)
*       88 = UAC85/U238/VDD (-1535.5 , 588)
*       88 = UAC85/U245/Vdd (-1480 , 588.5)
*       88 = UAC85/U218/VDD (-1456 , 585.5)
*       88 = UAC85/U235/VDD (-1309 , 588)
*       88 = UAC85/U229/Vdd (-1346 , 588.5)
*       88 = UAC85/U254/Vdd (-1416 , 544.5)
*       88 = UAC85/U253/VDD (-1330 , 542.5)
*       88 = UAC85/U247/Vdd (-1302 , 544.5)
*       88 = UAC85/U246/Vdd (-1254 , 544.5)
*       88 = UAC85/U236/VDD (-1264.5 , 588)
*       88 = UAC55/U262/VDD (-1127 , 633)
*       88 = UAC55/U219/VDD (-1163.5 , 632)
*       88 = UAC55/U222/VDD (-1091 , 629.5)
*       88 = UAC55/U220/VDD (-992 , 632)
*       88 = UAC55/U206/VDD (-960.5 , 629.5)
*       88 = UAC55/U246/Vdd (-882.5 , 544.5)
*       88 = UAC55/U254/Vdd (-1044.5 , 544.5)
*       88 = UAC55/U253/VDD (-958.5 , 542.5)
*       88 = UAC55/U247/Vdd (-930.5 , 544.5)
*       88 = UAC55/U245/Vdd (-1108.5 , 588.5)
*       88 = UAC55/U238/VDD (-1164 , 588)
*       88 = UAC55/U218/VDD (-1084.5 , 585.5)
*       88 = UAC55/U236/VDD (-893 , 588)
*       88 = UAC55/U235/VDD (-937.5 , 588)
*       88 = UAC55/U229/Vdd (-974.5 , 588.5)
*       88 = UAC56/U219/VDD (-800 , 632)
*       88 = UAC56/U262/VDD (-763.5 , 633)
*       88 = UAC56/U222/VDD (-727.5 , 629.5)
*       88 = UAC56/U206/VDD (-597 , 629.5)
*       88 = UAC56/U220/VDD (-628.5 , 632)
*       88 = UAC56/U254/Vdd (-681 , 544.5)
*       88 = UAC56/U253/VDD (-595 , 542.5)
*       88 = UAC56/U238/VDD (-800.5 , 588)
*       88 = UAC56/U245/Vdd (-745 , 588.5)
*       88 = UAC56/U218/VDD (-721 , 585.5)
*       88 = UAC56/U229/Vdd (-611 , 588.5)
*       88 = UAC56/U247/Vdd (-567 , 544.5)
*       88 = UAC56/U246/Vdd (-519 , 544.5)
*       88 = UAC56/U236/VDD (-529.5 , 588)
*       88 = UAC56/U235/VDD (-574 , 588)
*       88 = UAC57/U262/VDD (-399 , 633)
*       88 = UAC57/U219/VDD (-435.5 , 632)
*       88 = UAC57/U222/VDD (-363 , 629.5)
*       88 = UAC57/U206/VDD (-232.5 , 629.5)
*       88 = UAC57/U220/VDD (-264 , 632)
*       88 = UAC57/U238/VDD (-436 , 588)
*       88 = UAC57/U245/Vdd (-380.5 , 588.5)
*       88 = UAC57/U218/VDD (-356.5 , 585.5)
*       88 = UAC57/U235/VDD (-209.5 , 588)
*       88 = UAC57/U229/Vdd (-246.5 , 588.5)
*       88 = UAC57/U254/Vdd (-316.5 , 544.5)
*       88 = UAC57/U253/VDD (-230.5 , 542.5)
*       88 = UAC57/U247/Vdd (-202.5 , 544.5)
*       88 = UAC57/U246/Vdd (-154.5 , 544.5)
*       88 = UAC57/U236/VDD (-165 , 588)
*       88 = UAC58/U262/VDD (-35.5 , 633)
*       88 = UAC58/U222/VDD (0.5 , 629.5)
*       88 = UAC58/U219/VDD (-72 , 632)
*       88 = UAC58/U220/VDD (99.5 , 632)
*       88 = UAC58/U206/VDD (131 , 629.5)
*       88 = UAC54/U254/Vdd (47.5 , 707)
*       88 = UAC54/U253/VDD (133.5 , 705)
*       88 = UAC54/U247/Vdd (161.5 , 707)
*       88 = UAC58/U254/Vdd (47 , 544.5)
*       88 = UAC58/U253/VDD (133 , 542.5)
*       88 = UAC58/U247/Vdd (161 , 544.5)
*       88 = UAC58/U236/VDD (198.5 , 588)
*       88 = UAC58/U235/VDD (154 , 588)
*       88 = UAC58/U229/Vdd (117 , 588.5)
*       88 = UAC58/U245/Vdd (-17 , 588.5)
*       88 = UAC58/U238/VDD (-72.5 , 588)
*       88 = UAC58/U218/VDD (7 , 585.5)
*       88 = UAC61/U220/VDD (99 , 469.5)
*       88 = UAC60/U222/VDD (-363.5 , 467)
*       88 = UAC66/U236/VDD (-530 , 425.5)
*       88 = UAC66/U235/VDD (-574.5 , 425.5)
*       88 = UAC91/U222/VDD (-1463 , 467)
*       88 = UAC92/U236/VDD (-1633 , 425.5)
*       88 = UAC92/U235/VDD (-1677.5 , 425.5)
*       88 = UAC93/U222/VDD (-2191.002 , 467)
*       88 = UAC93/U220/VDD (-2096 , 469.5)
*       88 = UAC95/U236/VDD (-2734.5 , 425.5)
*       88 = UAC95/U235/VDD (-2779 , 425.5)
*       88 = UAC119/U231/VDD (-3393 , 379)
*       88 = UAC119/U224/Vdd (-3408 , 425)
*       88 = UAC119/U220/VDD (-3318 , 376.5)
*       88 = UAC119/U232/Vdd (-3345 , 380)
*       88 = UAC119/U226/Vdd (-3324 , 425)
*       88 = UAC119/U225/VDD (-3372 , 424)
*       88 = UAC119/U230/Vdd (-3240 , 425)
*       88 = UAC119/U229/VDD (-3288 , 424)
*       88 = UAC119/U222/VDD (-3401 , 469.5)
*       88 = UAC119/U223/Vdd (-3353 , 470.5)
*       88 = UAC119/U228/Vdd (-3261 , 470.5)
*       88 = UAC119/U227/VDD (-3279.5 , 468)
*       88 = UAC95/U219/VDD (-3005 , 469.5)
*       88 = UAC95/U262/VDD (-2968.5 , 470.5)
*       88 = UAC95/U222/VDD (-2932.5 , 467)
*       88 = UAC95/U206/VDD (-2802 , 467)
*       88 = UAC95/U220/VDD (-2833.5 , 469.5)
*       88 = UAC95/U247/Vdd (-2772 , 382)
*       88 = UAC95/U246/Vdd (-2724 , 382)
*       88 = UAC95/U254/Vdd (-2886 , 382)
*       88 = UAC95/U253/VDD (-2800 , 380)
*       88 = UAC95/U218/VDD (-2926 , 423)
*       88 = UAC95/U238/VDD (-3005.5 , 425.5)
*       88 = UAC95/U245/Vdd (-2950 , 426)
*       88 = UAC95/U229/Vdd (-2816 , 426)
*       88 = UAC94/U262/VDD (-2601.5 , 470.5)
*       88 = UAC94/U219/VDD (-2638 , 469.5)
*       88 = UAC94/U222/VDD (-2565.5 , 467)
*       88 = UAC94/U206/VDD (-2435 , 467)
*       88 = UAC94/U220/VDD (-2466.5 , 469.5)
*       88 = UAC94/U218/VDD (-2559 , 423)
*       88 = UAC94/U254/Vdd (-2519 , 382)
*       88 = UAC94/U253/VDD (-2433 , 380)
*       88 = UAC94/U247/Vdd (-2405 , 382)
*       88 = UAC94/U246/Vdd (-2357 , 382)
*       88 = UAC94/U238/VDD (-2638.5 , 425.5)
*       88 = UAC94/U245/Vdd (-2583 , 426)
*       88 = UAC94/U235/VDD (-2412 , 425.5)
*       88 = UAC94/U229/Vdd (-2449 , 426)
*       88 = UAC94/U236/VDD (-2367.5 , 425.5)
*       88 = UAC93/U262/VDD (-2231 , 470.5)
*       88 = UAC93/U219/VDD (-2267.5 , 469.5)
*       88 = UAC93/U206/VDD (-2064.5 , 467)
*       88 = UAC93/U254/Vdd (-2148.5 , 382)
*       88 = UAC93/U253/VDD (-2062.5 , 380)
*       88 = UAC93/U247/Vdd (-2034.5 , 382)
*       88 = UAC93/U218/VDD (-2188.5 , 423)
*       88 = UAC93/U246/Vdd (-1986.5 , 382)
*       88 = UAC93/U245/Vdd (-2212.5 , 426)
*       88 = UAC93/U238/VDD (-2268 , 425.5)
*       88 = UAC93/U236/VDD (-1997 , 425.5)
*       88 = UAC93/U235/VDD (-2041.5 , 425.5)
*       88 = UAC93/U229/Vdd (-2078.5 , 426)
*       88 = UAC92/U219/VDD (-1903.5 , 469.5)
*       88 = UAC92/U262/VDD (-1867 , 470.5)
*       88 = UAC92/U222/VDD (-1831 , 467)
*       88 = UAC92/U206/VDD (-1700.5 , 467)
*       88 = UAC92/U220/VDD (-1732 , 469.5)
*       88 = UAC92/U247/Vdd (-1670.5 , 382)
*       88 = UAC92/U246/Vdd (-1622.5 , 382)
*       88 = UAC92/U254/Vdd (-1784.5 , 382)
*       88 = UAC92/U253/VDD (-1698.5 , 380)
*       88 = UAC92/U218/VDD (-1824.5 , 423)
*       88 = UAC92/U238/VDD (-1904 , 425.5)
*       88 = UAC92/U245/Vdd (-1848.5 , 426)
*       88 = UAC92/U229/Vdd (-1714.5 , 426)
*       88 = UAC91/U262/VDD (-1499 , 470.5)
*       88 = UAC91/U219/VDD (-1535.5 , 469.5)
*       88 = UAC91/U206/VDD (-1332.5 , 467)
*       88 = UAC91/U220/VDD (-1364 , 469.5)
*       88 = UAC91/U218/VDD (-1456.5 , 423)
*       88 = UAC91/U254/Vdd (-1416.5 , 382)
*       88 = UAC91/U253/VDD (-1330.5 , 380)
*       88 = UAC91/U247/Vdd (-1302.5 , 382)
*       88 = UAC91/U246/Vdd (-1254.5 , 382)
*       88 = UAC91/U238/VDD (-1536 , 425.5)
*       88 = UAC91/U245/Vdd (-1480.5 , 426)
*       88 = UAC91/U235/VDD (-1309.5 , 425.5)
*       88 = UAC91/U229/Vdd (-1346.5 , 426)
*       88 = UAC91/U236/VDD (-1265 , 425.5)
*       88 = UAC59/U262/VDD (-1127.5 , 470.5)
*       88 = UAC59/U222/VDD (-1091.5 , 467)
*       88 = UAC59/U219/VDD (-1164 , 469.5)
*       88 = UAC59/U220/VDD (-992.5 , 469.5)
*       88 = UAC59/U206/VDD (-961 , 467)
*       88 = UAC59/U246/Vdd (-883 , 382)
*       88 = UAC59/U254/Vdd (-1045 , 382)
*       88 = UAC59/U253/VDD (-959 , 380)
*       88 = UAC59/U247/Vdd (-931 , 382)
*       88 = UAC59/U218/VDD (-1085 , 423)
*       88 = UAC59/U245/Vdd (-1109 , 426)
*       88 = UAC59/U238/VDD (-1164.5 , 425.5)
*       88 = UAC59/U236/VDD (-893.5 , 425.5)
*       88 = UAC59/U235/VDD (-938 , 425.5)
*       88 = UAC59/U229/Vdd (-975 , 426)
*       88 = UAC66/U219/VDD (-800.5 , 469.5)
*       88 = UAC66/U262/VDD (-764 , 470.5)
*       88 = UAC66/U222/VDD (-728 , 467)
*       88 = UAC66/U206/VDD (-597.5 , 467)
*       88 = UAC66/U220/VDD (-629 , 469.5)
*       88 = UAC66/U254/Vdd (-681.5 , 382)
*       88 = UAC66/U253/VDD (-595.5 , 380)
*       88 = UAC66/U218/VDD (-721.5 , 423)
*       88 = UAC66/U247/Vdd (-567.5 , 382)
*       88 = UAC66/U246/Vdd (-519.5 , 382)
*       88 = UAC66/U238/VDD (-801 , 425.5)
*       88 = UAC66/U245/Vdd (-745.5 , 426)
*       88 = UAC66/U229/Vdd (-611.5 , 426)
*       88 = UAC60/U262/VDD (-399.5 , 470.5)
*       88 = UAC60/U219/VDD (-436 , 469.5)
*       88 = UAC60/U206/VDD (-233 , 467)
*       88 = UAC60/U220/VDD (-264.5 , 469.5)
*       88 = UAC60/U218/VDD (-357 , 423)
*       88 = UAC60/U254/Vdd (-317 , 382)
*       88 = UAC60/U253/VDD (-231 , 380)
*       88 = UAC60/U247/Vdd (-203 , 382)
*       88 = UAC60/U246/Vdd (-155 , 382)
*       88 = UAC60/U238/VDD (-436.5 , 425.5)
*       88 = UAC60/U245/Vdd (-381 , 426)
*       88 = UAC60/U235/VDD (-210 , 425.5)
*       88 = UAC60/U229/Vdd (-247 , 426)
*       88 = UAC60/U236/VDD (-165.5 , 425.5)
*       88 = UAC61/U262/VDD (-36 , 470.5)
*       88 = UAC61/U222/VDD (0 , 467)
*       88 = UAC61/U219/VDD (-72.5 , 469.5)
*       88 = UAC61/U206/VDD (130.5 , 467)
*       88 = UAC61/U254/Vdd (46.5 , 382)
*       88 = UAC61/U253/VDD (132.5 , 380)
*       88 = UAC61/U247/Vdd (160.5 , 382)
*       88 = UAC61/U246/Vdd (208.5 , 382)
*       88 = UAC61/U218/VDD (6.5 , 423)
*       88 = UAC65/U245/Vdd (-18 , 263.5)
*       88 = UAC65/U238/VDD (-73.5 , 263)
*       88 = UAC65/U218/VDD (6 , 260.5)
*       88 = UAC65/U236/VDD (197.5 , 263)
*       88 = UAC65/U235/VDD (153 , 263)
*       88 = UAC65/U229/Vdd (116 , 263.5)
*       88 = UAC65/U220/VDD (98.5 , 307)
*       88 = UAC64/U238/VDD (-437 , 263)
*       88 = UAC64/U245/Vdd (-381.5 , 263.5)
*       88 = UAC64/U218/VDD (-357.5 , 260.5)
*       88 = UAC64/U235/VDD (-210.5 , 263)
*       88 = UAC64/U229/Vdd (-247.5 , 263.5)
*       88 = UAC64/U222/VDD (-364 , 304.5)
*       88 = UAC63/U236/VDD (-530.5 , 263)
*       88 = UAC63/U235/VDD (-575 , 263)
*       88 = UAC63/U238/VDD (-801.5 , 263)
*       88 = UAC63/U245/Vdd (-746 , 263.5)
*       88 = UAC63/U218/VDD (-722 , 260.5)
*       88 = UAC63/U229/Vdd (-612 , 263.5)
*       88 = UAC62/U245/Vdd (-1109.5 , 263.5)
*       88 = UAC62/U238/VDD (-1165 , 263)
*       88 = UAC62/U218/VDD (-1085.5 , 260.5)
*       88 = UAC62/U236/VDD (-894 , 263)
*       88 = UAC62/U235/VDD (-938.5 , 263)
*       88 = UAC62/U229/Vdd (-975.5 , 263.5)
*       88 = UAC96/U238/VDD (-1536.5 , 263)
*       88 = UAC96/U245/Vdd (-1481 , 263.5)
*       88 = UAC96/U218/VDD (-1457 , 260.5)
*       88 = UAC96/U235/VDD (-1310 , 263)
*       88 = UAC96/U229/Vdd (-1347 , 263.5)
*       88 = UAC96/U222/VDD (-1463.5 , 304.5)
*       88 = UAC97/U236/VDD (-1633.5 , 263)
*       88 = UAC97/U235/VDD (-1678 , 263)
*       88 = UAC97/U238/VDD (-1904.5 , 263)
*       88 = UAC97/U245/Vdd (-1849 , 263.5)
*       88 = UAC97/U218/VDD (-1825 , 260.5)
*       88 = UAC97/U229/Vdd (-1715 , 263.5)
*       88 = UAC98/U245/Vdd (-2213 , 263.5)
*       88 = UAC98/U238/VDD (-2268.5 , 263)
*       88 = UAC98/U218/VDD (-2189 , 260.5)
*       88 = UAC98/U236/VDD (-1997.5 , 263)
*       88 = UAC98/U235/VDD (-2042 , 263)
*       88 = UAC98/U229/Vdd (-2079 , 263.5)
*       88 = UAC98/U222/VDD (-2191.002 , 304.5)
*       88 = UAC98/U220/VDD (-2096.5 , 307)
*       88 = UAC99/U245/Vdd (-2583.5 , 263.5)
*       88 = UAC99/U218/VDD (-2559.5 , 260.5)
*       88 = UAC99/U238/VDD (-2639 , 263)
*       88 = UAC99/U235/VDD (-2412.5 , 263)
*       88 = UAC99/U229/Vdd (-2449.5 , 263.5)
*       88 = UAC100/U236/VDD (-2735 , 263)
*       88 = UAC100/U235/VDD (-2779.5 , 263)
*       88 = UAC100/U238/VDD (-3006 , 263)
*       88 = UAC100/U245/Vdd (-2950.5 , 263.5)
*       88 = UAC100/U218/VDD (-2926.5 , 260.5)
*       88 = UAC100/U229/Vdd (-2816.5 , 263.5)
*       88 = UAC101/U245/Vdd (-3322 , 263.5)
*       88 = UAC101/U238/VDD (-3377.5 , 263)
*       88 = UAC101/U218/VDD (-3298 , 260.5)
*       88 = UAC101/U236/VDD (-3106.5 , 263)
*       88 = UAC101/U235/VDD (-3151 , 263)
*       88 = UAC101/U229/Vdd (-3188 , 263.5)
*       88 = UAC101/U220/VDD (-3205.5 , 307)
*       88 = UAC120/U232/Vdd (-3710 , 217.5)
*       88 = UAC120/U231/VDD (-3758 , 216.5)
*       88 = UAC120/U220/VDD (-3683 , 214)
*       88 = UAC120/U225/VDD (-3737 , 261.5)
*       88 = UAC120/U224/Vdd (-3773 , 262.5)
*       88 = UAC120/U223/Vdd (-3718 , 308)
*       88 = UAC120/U222/VDD (-3766 , 307)
*       88 = UAC120/U230/Vdd (-3605 , 262.5)
*       88 = UAC120/U229/VDD (-3653 , 261.5)
*       88 = UAC120/U226/Vdd (-3689 , 262.5)
*       88 = UAC120/U228/Vdd (-3626 , 308)
*       88 = UAC120/U227/VDD (-3644.5 , 305.5)
*       88 = UAC101/U262/VDD (-3340.5 , 308)
*       88 = UAC101/U222/VDD (-3304.5 , 304.5)
*       88 = UAC101/U219/VDD (-3377 , 307)
*       88 = UAC101/U206/VDD (-3174 , 304.5)
*       88 = UAC101/U254/Vdd (-3258 , 219.5)
*       88 = UAC101/U253/VDD (-3172 , 217.5)
*       88 = UAC101/U247/Vdd (-3144 , 219.5)
*       88 = UAC101/U246/Vdd (-3096 , 219.5)
*       88 = UAC100/U219/VDD (-3005.5 , 307)
*       88 = UAC100/U262/VDD (-2969 , 308)
*       88 = UAC100/U222/VDD (-2933 , 304.5)
*       88 = UAC100/U206/VDD (-2802.5 , 304.5)
*       88 = UAC100/U220/VDD (-2834 , 307)
*       88 = UAC100/U247/Vdd (-2772.5 , 219.5)
*       88 = UAC100/U246/Vdd (-2724.5 , 219.5)
*       88 = UAC100/U254/Vdd (-2886.5 , 219.5)
*       88 = UAC100/U253/VDD (-2800.5 , 217.5)
*       88 = UAC99/U262/VDD (-2602 , 308)
*       88 = UAC99/U219/VDD (-2638.5 , 307)
*       88 = UAC99/U222/VDD (-2566 , 304.5)
*       88 = UAC99/U206/VDD (-2435.5 , 304.5)
*       88 = UAC99/U220/VDD (-2467 , 307)
*       88 = UAC99/U254/Vdd (-2519.5 , 219.5)
*       88 = UAC99/U253/VDD (-2433.5 , 217.5)
*       88 = UAC99/U247/Vdd (-2405.5 , 219.5)
*       88 = UAC99/U246/Vdd (-2357.5 , 219.5)
*       88 = UAC99/U236/VDD (-2368 , 263)
*       88 = UAC98/U262/VDD (-2231.5 , 308)
*       88 = UAC98/U219/VDD (-2268 , 307)
*       88 = UAC98/U206/VDD (-2065 , 304.5)
*       88 = UAC98/U254/Vdd (-2149 , 219.5)
*       88 = UAC98/U253/VDD (-2063 , 217.5)
*       88 = UAC98/U247/Vdd (-2035 , 219.5)
*       88 = UAC98/U246/Vdd (-1987 , 219.5)
*       88 = UAC97/U219/VDD (-1904 , 307)
*       88 = UAC97/U262/VDD (-1867.5 , 308)
*       88 = UAC97/U222/VDD (-1831.5 , 304.5)
*       88 = UAC97/U206/VDD (-1701 , 304.5)
*       88 = UAC97/U220/VDD (-1732.5 , 307)
*       88 = UAC97/U247/Vdd (-1671 , 219.5)
*       88 = UAC97/U246/Vdd (-1623 , 219.5)
*       88 = UAC97/U254/Vdd (-1785 , 219.5)
*       88 = UAC97/U253/VDD (-1699 , 217.5)
*       88 = UAC96/U262/VDD (-1499.5 , 308)
*       88 = UAC96/U219/VDD (-1536 , 307)
*       88 = UAC96/U206/VDD (-1333 , 304.5)
*       88 = UAC96/U220/VDD (-1364.5 , 307)
*       88 = UAC96/U254/Vdd (-1417 , 219.5)
*       88 = UAC96/U253/VDD (-1331 , 217.5)
*       88 = UAC96/U247/Vdd (-1303 , 219.5)
*       88 = UAC96/U246/Vdd (-1255 , 219.5)
*       88 = UAC96/U236/VDD (-1265.5 , 263)
*       88 = UAC62/U262/VDD (-1128 , 308)
*       88 = UAC62/U222/VDD (-1092 , 304.5)
*       88 = UAC62/U219/VDD (-1164.5 , 307)
*       88 = UAC62/U220/VDD (-993 , 307)
*       88 = UAC62/U206/VDD (-961.5 , 304.5)
*       88 = UAC62/U246/Vdd (-883.5 , 219.5)
*       88 = UAC62/U254/Vdd (-1045.5 , 219.5)
*       88 = UAC62/U253/VDD (-959.5 , 217.5)
*       88 = UAC62/U247/Vdd (-931.5 , 219.5)
*       88 = UAC63/U219/VDD (-801 , 307)
*       88 = UAC63/U262/VDD (-764.5 , 308)
*       88 = UAC63/U222/VDD (-728.5 , 304.5)
*       88 = UAC63/U206/VDD (-598 , 304.5)
*       88 = UAC63/U220/VDD (-629.5 , 307)
*       88 = UAC63/U254/Vdd (-682 , 219.5)
*       88 = UAC63/U253/VDD (-596 , 217.5)
*       88 = UAC63/U247/Vdd (-568 , 219.5)
*       88 = UAC63/U246/Vdd (-520 , 219.5)
*       88 = UAC64/U262/VDD (-400 , 308)
*       88 = UAC64/U219/VDD (-436.5 , 307)
*       88 = UAC64/U206/VDD (-233.5 , 304.5)
*       88 = UAC64/U220/VDD (-265 , 307)
*       88 = UAC64/U254/Vdd (-317.5 , 219.5)
*       88 = UAC64/U253/VDD (-231.5 , 217.5)
*       88 = UAC64/U247/Vdd (-203.5 , 219.5)
*       88 = UAC64/U246/Vdd (-155.5 , 219.5)
*       88 = UAC64/U236/VDD (-166 , 263)
*       88 = UAC65/U262/VDD (-36.5 , 308)
*       88 = UAC65/U222/VDD (-0.5 , 304.5)
*       88 = UAC65/U219/VDD (-73 , 307)
*       88 = UAC65/U206/VDD (130 , 304.5)
*       88 = UAC70/U220/VDD (98 , 145.5)
*       88 = UAC69/U222/VDD (-364.5 , 143)
*       88 = UAC102/U222/VDD (-1457.5 , 143)
*       88 = UAC103/U206/VDD (-1691.002 , 143)
*       88 = UAC104/U206/VDD (-2059 , 143)
*       88 = UAC104/U220/VDD (-2090.5 , 145.5)
*       88 = UAC105/U222/VDD (-2560 , 143)
*       88 = UAC106/U206/VDD (-2791.002 , 143)
*       88 = UAC107/U220/VDD (-3199.5 , 145.5)
*       88 = UAC121/U220/VDD (-3994 , 52.5)
*       88 = UAC121/U232/Vdd (-4021 , 56)
*       88 = UAC121/U231/VDD (-4069 , 55)
*       88 = UAC121/U226/Vdd (-4000 , 101)
*       88 = UAC121/U225/VDD (-4048 , 100)
*       88 = UAC121/U224/Vdd (-4084 , 101)
*       88 = UAC121/U230/Vdd (-3916 , 101)
*       88 = UAC121/U229/VDD (-3964 , 100)
*       88 = UAC121/U223/Vdd (-4029 , 146.5)
*       88 = UAC121/U222/VDD (-4077 , 145.5)
*       88 = UAC121/U228/Vdd (-3937 , 146.5)
*       88 = UAC121/U227/VDD (-3955.5 , 144)
*       88 = UAC109/U262/VDD (-3707 , 146.5)
*       88 = UAC109/U219/VDD (-3743.5 , 145.5)
*       88 = UAC109/U222/VDD (-3671 , 143)
*       88 = UAC109/U206/VDD (-3540.5 , 143)
*       88 = UAC109/U220/VDD (-3572 , 145.5)
*       88 = UAC109/U253/VDD (-3538.5 , 56)
*       88 = UAC109/U247/Vdd (-3510.5 , 58)
*       88 = UAC109/U254/Vdd (-3624.5 , 58)
*       88 = UAC109/U238/VDD (-3744 , 101.5)
*       88 = UAC109/U245/Vdd (-3688.5 , 102)
*       88 = UAC109/U218/VDD (-3664.5 , 99)
*       88 = UAC109/U235/VDD (-3517.5 , 101.5)
*       88 = UAC109/U229/Vdd (-3554.5 , 102)
*       88 = UAC109/U246/Vdd (-3462.5 , 58)
*       88 = UAC109/U236/VDD (-3473 , 101.5)
*       88 = UAC107/U262/VDD (-3334.5 , 146.5)
*       88 = UAC107/U222/VDD (-3298.5 , 143)
*       88 = UAC107/U219/VDD (-3371 , 145.5)
*       88 = UAC107/U206/VDD (-3168 , 143)
*       88 = UAC107/U254/Vdd (-3252 , 58)
*       88 = UAC107/U253/VDD (-3166 , 56)
*       88 = UAC107/U247/Vdd (-3138 , 58)
*       88 = UAC107/U245/Vdd (-3316 , 102)
*       88 = UAC107/U238/VDD (-3371.5 , 101.5)
*       88 = UAC107/U218/VDD (-3292 , 99)
*       88 = UAC107/U236/VDD (-3100.5 , 101.5)
*       88 = UAC107/U235/VDD (-3145 , 101.5)
*       88 = UAC107/U229/Vdd (-3182 , 102)
*       88 = UAC107/U246/Vdd (-3090 , 58)
*       88 = UAC106/U219/VDD (-2999.5 , 145.5)
*       88 = UAC106/U262/VDD (-2963 , 146.5)
*       88 = UAC106/U222/VDD (-2927 , 143)
*       88 = UAC106/U220/VDD (-2828 , 145.5)
*       88 = UAC106/U254/Vdd (-2880.5 , 58)
*       88 = UAC106/U253/VDD (-2794.5 , 56)
*       88 = UAC106/U238/VDD (-3000 , 101.5)
*       88 = UAC106/U245/Vdd (-2944.5 , 102)
*       88 = UAC106/U218/VDD (-2920.5 , 99)
*       88 = UAC106/U229/Vdd (-2810.5 , 102)
*       88 = UAC106/U247/Vdd (-2766.5 , 58)
*       88 = UAC106/U246/Vdd (-2718.5 , 58)
*       88 = UAC106/U236/VDD (-2729 , 101.5)
*       88 = UAC106/U235/VDD (-2773.5 , 101.5)
*       88 = UAC105/U262/VDD (-2596 , 146.5)
*       88 = UAC105/U219/VDD (-2632.5 , 145.5)
*       88 = UAC105/U206/VDD (-2429.5 , 143)
*       88 = UAC105/U220/VDD (-2461 , 145.5)
*       88 = UAC105/U238/VDD (-2633 , 101.5)
*       88 = UAC105/U245/Vdd (-2577.5 , 102)
*       88 = UAC105/U218/VDD (-2553.5 , 99)
*       88 = UAC105/U235/VDD (-2406.5 , 101.5)
*       88 = UAC105/U229/Vdd (-2443.5 , 102)
*       88 = UAC105/U254/Vdd (-2513.5 , 58)
*       88 = UAC105/U253/VDD (-2427.5 , 56)
*       88 = UAC105/U247/Vdd (-2399.5 , 58)
*       88 = UAC105/U246/Vdd (-2351.5 , 58)
*       88 = UAC105/U236/VDD (-2362 , 101.5)
*       88 = UAC104/U262/VDD (-2225.5 , 146.5)
*       88 = UAC104/U219/VDD (-2262 , 145.5)
*       88 = UAC104/U222/VDD (-2189.5 , 143)
*       88 = UAC104/U246/Vdd (-1981 , 58)
*       88 = UAC104/U254/Vdd (-2143 , 58)
*       88 = UAC104/U253/VDD (-2057 , 56)
*       88 = UAC104/U247/Vdd (-2029 , 58)
*       88 = UAC104/U236/VDD (-1991.5 , 101.5)
*       88 = UAC104/U235/VDD (-2036 , 101.5)
*       88 = UAC104/U229/Vdd (-2073 , 102)
*       88 = UAC104/U245/Vdd (-2207 , 102)
*       88 = UAC104/U238/VDD (-2262.5 , 101.5)
*       88 = UAC104/U218/VDD (-2183 , 99)
*       88 = UAC103/U219/VDD (-1898 , 145.5)
*       88 = UAC103/U262/VDD (-1861.5 , 146.5)
*       88 = UAC103/U222/VDD (-1825.5 , 143)
*       88 = UAC103/U220/VDD (-1726.5 , 145.5)
*       88 = UAC103/U254/Vdd (-1779 , 58)
*       88 = UAC103/U253/VDD (-1693 , 56)
*       88 = UAC103/U247/Vdd (-1665 , 58)
*       88 = UAC103/U246/Vdd (-1617 , 58)
*       88 = UAC103/U238/VDD (-1898.5 , 101.5)
*       88 = UAC103/U245/Vdd (-1843 , 102)
*       88 = UAC103/U218/VDD (-1819 , 99)
*       88 = UAC103/U229/Vdd (-1709 , 102)
*       88 = UAC103/U236/VDD (-1627.5 , 101.5)
*       88 = UAC103/U235/VDD (-1672 , 101.5)
*       88 = UAC102/U262/VDD (-1493.5 , 146.5)
*       88 = UAC102/U219/VDD (-1530 , 145.5)
*       88 = UAC102/U206/VDD (-1327 , 143)
*       88 = UAC102/U220/VDD (-1358.5 , 145.5)
*       88 = UAC102/U238/VDD (-1530.5 , 101.5)
*       88 = UAC102/U245/Vdd (-1475 , 102)
*       88 = UAC102/U218/VDD (-1451 , 99)
*       88 = UAC102/U235/VDD (-1304 , 101.5)
*       88 = UAC102/U229/Vdd (-1341 , 102)
*       88 = UAC102/U254/Vdd (-1411 , 58)
*       88 = UAC102/U253/VDD (-1325 , 56)
*       88 = UAC102/U247/Vdd (-1297 , 58)
*       88 = UAC102/U246/Vdd (-1249 , 58)
*       88 = UAC102/U236/VDD (-1259.5 , 101.5)
*       88 = UAC67/U262/VDD (-1128.5 , 146.5)
*       88 = UAC67/U222/VDD (-1092.5 , 143)
*       88 = UAC67/U219/VDD (-1165 , 145.5)
*       88 = UAC67/U220/VDD (-993.5 , 145.5)
*       88 = UAC67/U206/VDD (-962 , 143)
*       88 = UAC67/U254/Vdd (-1046 , 58)
*       88 = UAC67/U253/VDD (-960 , 56)
*       88 = UAC67/U247/Vdd (-932 , 58)
*       88 = UAC67/U245/Vdd (-1110 , 102)
*       88 = UAC67/U238/VDD (-1165.5 , 101.5)
*       88 = UAC67/U218/VDD (-1086 , 99)
*       88 = UAC67/U236/VDD (-894.5 , 101.5)
*       88 = UAC67/U235/VDD (-939 , 101.5)
*       88 = UAC67/U229/Vdd (-976 , 102)
*       88 = UAC67/U246/Vdd (-884 , 58)
*       88 = UAC68/U219/VDD (-801.5 , 145.5)
*       88 = UAC68/U262/VDD (-765 , 146.5)
*       88 = UAC68/U222/VDD (-729 , 143)
*       88 = UAC68/U206/VDD (-598.5 , 143)
*       88 = UAC68/U220/VDD (-630 , 145.5)
*       88 = UAC68/U254/Vdd (-682.5 , 58)
*       88 = UAC68/U253/VDD (-596.5 , 56)
*       88 = UAC68/U238/VDD (-802 , 101.5)
*       88 = UAC68/U245/Vdd (-746.5 , 102)
*       88 = UAC68/U218/VDD (-722.5 , 99)
*       88 = UAC68/U229/Vdd (-612.5 , 102)
*       88 = UAC68/U247/Vdd (-568.5 , 58)
*       88 = UAC68/U246/Vdd (-520.5 , 58)
*       88 = UAC68/U236/VDD (-531 , 101.5)
*       88 = UAC68/U235/VDD (-575.5 , 101.5)
*       88 = UAC69/U262/VDD (-400.5 , 146.5)
*       88 = UAC69/U219/VDD (-437 , 145.5)
*       88 = UAC69/U206/VDD (-234 , 143)
*       88 = UAC69/U220/VDD (-265.5 , 145.5)
*       88 = UAC69/U238/VDD (-437.5 , 101.5)
*       88 = UAC69/U245/Vdd (-382 , 102)
*       88 = UAC69/U218/VDD (-358 , 99)
*       88 = UAC69/U235/VDD (-211 , 101.5)
*       88 = UAC69/U229/Vdd (-248 , 102)
*       88 = UAC69/U254/Vdd (-318 , 58)
*       88 = UAC69/U253/VDD (-232 , 56)
*       88 = UAC69/U247/Vdd (-204 , 58)
*       88 = UAC69/U246/Vdd (-156 , 58)
*       88 = UAC69/U236/VDD (-166.5 , 101.5)
*       88 = UAC70/U262/VDD (-37 , 146.5)
*       88 = UAC70/U222/VDD (-1 , 143)
*       88 = UAC70/U219/VDD (-73.5 , 145.5)
*       88 = UAC70/U206/VDD (129.5 , 143)
*       88 = UAC65/U254/Vdd (46 , 219.5)
*       88 = UAC65/U253/VDD (132 , 217.5)
*       88 = UAC65/U247/Vdd (160 , 219.5)
*       88 = UAC65/U246/Vdd (208 , 219.5)
*       88 = UAC70/U218/VDD (8.997 , 99)
*       88 = UAC70/U245/Vdd (-18.5 , 102)
*       88 = UAC70/U238/VDD (-74 , 101.5)
*       88 = UAC70/U236/VDD (197 , 101.5)
*       88 = UAC70/U235/VDD (152.5 , 101.5)
*       88 = UAC70/U229/Vdd (115.5 , 102)
*       88 = UAC70/U254/Vdd (45.5 , 58)
*       88 = UAC70/U253/VDD (131.5 , 56)
*       88 = UAC70/U247/Vdd (159.5 , 58)
*       88 = UAC70/U246/Vdd (207.5 , 58)
*       88 = UAC74/U236/VDD (196.5 , -61)
*       88 = UAC74/U235/VDD (152 , -61)
*       88 = UAC74/U229/Vdd (115 , -60.5)
*       88 = UAC74/U245/Vdd (-19 , -60.5)
*       88 = UAC74/U238/VDD (-74.5 , -61)
*       88 = UAC74/U218/VDD (5 , -63.5)
*       88 = UAC74/U220/VDD (97.5 , -17)
*       88 = UAC73/U245/Vdd (-382.5 , -60.5)
*       88 = UAC73/U218/VDD (-358.5 , -63.5)
*       88 = UAC73/U238/VDD (-438 , -61)
*       88 = UAC73/U235/VDD (-211.5 , -61)
*       88 = UAC73/U229/Vdd (-248.5 , -60.5)
*       88 = UAC73/U222/VDD (-365 , -19.5)
*       88 = UAC72/U236/VDD (-531.5 , -61)
*       88 = UAC72/U235/VDD (-576 , -61)
*       88 = UAC72/U238/VDD (-802.5 , -61)
*       88 = UAC72/U245/Vdd (-747 , -60.5)
*       88 = UAC72/U218/VDD (-723 , -63.5)
*       88 = UAC72/U229/Vdd (-613 , -60.5)
*       88 = UAC71/U236/VDD (-895 , -61)
*       88 = UAC71/U235/VDD (-939.5 , -61)
*       88 = UAC71/U229/Vdd (-976.5 , -60.5)
*       88 = UAC71/U245/Vdd (-1110.5 , -60.5)
*       88 = UAC71/U238/VDD (-1166 , -61)
*       88 = UAC71/U218/VDD (-1086.5 , -63.5)
*       88 = UAC126/Vdd (-1340 , -16.5)
*       88 = UAC125/VDD (-1301.5 , -17)
*       88 = UAC124/Vdd (-1246 , -16.5)
*       88 = UAC71/U262/VDD (-1129 , -16)
*       88 = UAC71/U222/VDD (-1093 , -19.5)
*       88 = UAC71/U219/VDD (-1165.5 , -17)
*       88 = UAC71/U220/VDD (-994 , -17)
*       88 = UAC71/U206/VDD (-962.5 , -19.5)
*       88 = UAC72/U219/VDD (-802 , -17)
*       88 = UAC71/U254/Vdd (-1046.5 , -104.5)
*       88 = UAC71/U253/VDD (-960.5 , -106.5)
*       88 = UAC71/U247/Vdd (-932.5 , -104.5)
*       88 = UAC71/U246/Vdd (-884.5 , -104.5)
*       88 = UAC72/U262/VDD (-765.5 , -16)
*       88 = UAC72/U222/VDD (-729.5 , -19.5)
*       88 = UAC72/U206/VDD (-599 , -19.5)
*       88 = UAC72/U220/VDD (-630.5 , -17)
*       88 = UAC72/U254/Vdd (-683 , -104.5)
*       88 = UAC72/U253/VDD (-597 , -106.5)
*       88 = UAC72/U247/Vdd (-569 , -104.5)
*       88 = UAC72/U246/Vdd (-521 , -104.5)
*       88 = UAC73/U262/VDD (-401 , -16)
*       88 = UAC73/U219/VDD (-437.5 , -17)
*       88 = UAC73/U206/VDD (-234.5 , -19.5)
*       88 = UAC73/U220/VDD (-266 , -17)
*       88 = UAC73/U236/VDD (-167 , -61)
*       88 = UAC73/U254/Vdd (-318.5 , -104.5)
*       88 = UAC73/U253/VDD (-232.5 , -106.5)
*       88 = UAC73/U247/Vdd (-204.5 , -104.5)
*       88 = UAC73/U246/Vdd (-156.5 , -104.5)
*       88 = UAC74/U262/VDD (-37.5 , -16)
*       88 = UAC74/U222/VDD (-1.5 , -19.5)
*       88 = UAC74/U219/VDD (-74 , -17)
*       88 = UAC74/U206/VDD (129 , -19.5)
*       88 = UAC74/U254/Vdd (45 , -104.5)
*       88 = UAC74/U253/VDD (131 , -106.5)
*       88 = UAC74/U247/Vdd (159 , -104.5)
*       88 = UAC74/U246/Vdd (207 , -104.5)
*       88 = UAC61/U245/Vdd (-17.5 , 426)
*       88 = UAC61/U238/VDD (-73 , 425.5)
*       88 = UAC61/U236/VDD (198 , 425.5)
*       88 = UAC61/U235/VDD (153.5 , 425.5)
*       88 = UAC61/U229/Vdd (116.5 , 426)
*       88 = UAC58/U246/Vdd (209 , 544.5)
*       88 = UAC54/U246/Vdd (209.5 , 707)
*       88 = UAC42/U246/Vdd (210 , 868.5)
*       88 = UAC38/U254/Vdd (48.5 , 1031)
*       88 = UAC38/U253/VDD (134.5 , 1029)
*       88 = UAC38/U247/Vdd (162.5 , 1031)
*       88 = UAC38/U246/Vdd (210.5 , 1031)
*       88 = UAC34/U246/Vdd (211 , 1193.5)
*       94 = UAC34/U218/B (86 , 1215.5)
*       94 = UAC34/U229/Vout (125 , 1217)
*       95 = UAC34/U253/B (97.5 , 1162)
*       95 = UAC34/U246/Vout (217 , 1173)
*       96 = UAC34/U218/A (12.5 , 1220.5)
*       96 = UAC34/U222/Vout (41.5 , 1271.5)
*       98 = UAC34/U254/Vin (41 , 1173)
*       98 = UAC34/U253/OUT (75.5 , 1161.5)
*       101 = UAC34/U245/Vout (-9 , 1217)
*       101 = UAC34/U253/A (85 , 1161.5)
*       102 = UAC34/U245/Vin (-23 , 1217)
*       102 = UAC34/U238/OUT (-62.5 , 1204)
*       103 = UAC42/U219/A (-76.5 , 934.5)
*       103 = UAC38/B6 (-76.5 , 1024)
*       103 = UAC74/U238/A (-80 , -82.5)
*       103 = UAC74/B6 (-80 , -111.5)
*       103 = UAC74/U219/A (-79.5 , -38.5)
*       103 = UAC74/U235/A (146.5 , -82.5)
*       103 = UAC70/U238/A (-79.5 , 80)
*       103 = UAC70/U219/A (-79 , 124)
*       103 = UAC70/B6 (-79.5 , 51)
*       103 = UAC70/U235/A (147 , 80)
*       103 = UAC65/B6 (-79 , 212.5)
*       103 = UAC65/U238/A (-79 , 241.5)
*       103 = UAC65/U219/A (-78.5 , 285.5)
*       103 = UAC65/U235/A (147.5 , 241.5)
*       103 = UAC61/U238/A (-78.5 , 404)
*       103 = UAC61/B6 (-78.5 , 375)
*       103 = UAC61/U235/A (148 , 404)
*       103 = UAC61/U219/A (-78 , 448)
*       103 = UAC58/U238/A (-78 , 566.5)
*       103 = UAC58/U219/A (-77.5 , 610.5)
*       103 = UAC58/B6 (-78 , 537.5)
*       103 = UAC58/U235/A (148.5 , 566.5)
*       103 = UAC54/B6 (-77.5 , 700)
*       103 = UAC54/U238/A (-77.5 , 729)
*       103 = UAC54/U219/A (-77 , 773)
*       103 = UAC54/U235/A (149 , 729)
*       103 = UAC42/U238/A (-77 , 890.5)
*       103 = UAC42/B6 (-77 , 861.5)
*       103 = UAC42/U235/A (149.5 , 890.5)
*       103 = UAC38/U238/A (-76.5 , 1053)
*       103 = UAC38/U219/A (-76 , 1097)
*       103 = UAC38/U235/A (150 , 1053)
*       103 = UAC34/U238/A (-76 , 1215.5)
*       103 = UAC34/B6 (-76 , 1186.5)
*       103 = UAC34/U219/A (-75.5 , 1259.5)
*       103 = Bf0 (-75.5 , 1299)
*       103 = UAC34/U235/A (150.5 , 1215.5)
*       104 = UAC34/U238/B (-49.5 , 1215.5)
*       104 = UAC34/U220/A (96 , 1259.5)
*       104 = UAC34/C6 (96 , 1291.5)
*       104 = UAC32/U222/B (-648.5 , 1259.5)
*       104 = UAC32/U206/A (-591.5 , 1264.5)
*       104 = UAC31/U222/B (-1012 , 1259.5)
*       104 = UAC38/U238/B (-50 , 1053)
*       104 = UAC38/U220/A (95.5 , 1097)
*       104 = UAC79/U219/A (-1532 , 934.5)
*       104 = UAC78/B6 (-1532 , 1024)
*       104 = UAC102/U238/A (-1536 , 80)
*       104 = UAC102/U219/A (-1535.5 , 124)
*       104 = UAC102/B6 (-1536 , 51)
*       104 = UAC102/U235/A (-1309.5 , 80)
*       104 = UAC96/B6 (-1542 , 212.5)
*       104 = UAC96/U238/A (-1542 , 241.5)
*       104 = UAC96/U219/A (-1541.5 , 285.5)
*       104 = UAC96/U235/A (-1315.5 , 241.5)
*       104 = UAC91/U238/A (-1541.5 , 404)
*       104 = UAC91/B6 (-1541.5 , 375)
*       104 = UAC91/U235/A (-1315 , 404)
*       104 = UAC91/U219/A (-1541 , 448)
*       104 = UAC85/U238/A (-1541 , 566.5)
*       104 = UAC85/U219/A (-1540.5 , 610.5)
*       104 = UAC85/B6 (-1541 , 537.5)
*       104 = UAC85/U235/A (-1314.5 , 566.5)
*       104 = UAC81/B6 (-1540.5 , 700)
*       104 = UAC81/U238/A (-1540.5 , 729)
*       104 = UAC81/U219/A (-1540 , 773)
*       104 = UAC81/U235/A (-1314 , 729)
*       104 = UAC79/U238/A (-1532.5 , 890.5)
*       104 = UAC79/B6 (-1532.5 , 861.5)
*       104 = UAC79/U235/A (-1306 , 890.5)
*       104 = UAC42/U238/B (-50.5 , 890.5)
*       104 = UAC42/U220/A (95 , 934.5)
*       104 = UAC42/C6 (95 , 966.5)
*       104 = UAC42/U262/GND (-20.5 , 922)
*       104 = UAC42/U222/Gnd (1.5 , 919.5)
*       104 = UAC42/U219/GND (-41.5 , 922)
*       104 = UAC40/U262/GND (-748.5 , 922)
*       104 = UAC40/U222/Gnd (-726.5 , 919.5)
*       104 = UAC40/U219/GND (-769.5 , 922)
*       104 = UAC114/U223/GND (-2243 , 922.5)
*       104 = UAC114/U222/GND (-2260 , 922)
*       104 = UAC114/U224/GND (-2298 , 877)
*       104 = UAC54/U238/B (-51 , 729)
*       104 = UAC54/U220/A (94.5 , 773)
*       104 = UAC54/C6 (94.5 , 805)
*       104 = UAC54/U235/GND (184 , 716.5)
*       104 = UAC54/U229/Gnd (114.5 , 717)
*       104 = UAC54/U253/GND (133 , 674)
*       104 = UAC54/U247/Gnd (158.5 , 673)
*       104 = UAC54/U246/Gnd (206.5 , 673)
*       104 = UAC104/U238/A (-2268 , 80)
*       104 = UAC104/U219/A (-2267.5 , 124)
*       104 = UAC104/B6 (-2268 , 51)
*       104 = UAC104/U235/A (-2041.5 , 80)
*       104 = UAC98/B6 (-2274 , 212.5)
*       104 = UAC98/U238/A (-2274 , 241.5)
*       104 = UAC98/U219/A (-2273.5 , 285.5)
*       104 = UAC98/U235/A (-2047.5 , 241.5)
*       104 = UAC93/U238/A (-2273.5 , 404)
*       104 = UAC93/B6 (-2273.5 , 375)
*       104 = UAC93/U235/A (-2047 , 404)
*       104 = UAC93/U219/A (-2273 , 448)
*       104 = UAC88/U238/A (-2273 , 566.5)
*       104 = UAC88/U219/A (-2272.5 , 610.5)
*       104 = UAC88/B6 (-2273 , 537.5)
*       104 = UAC88/U235/A (-2046.5 , 566.5)
*       104 = UAC116/U230/GND (-2501 , 715.5)
*       104 = UAC116/U229/GND (-2518 , 715)
*       104 = UAC116/U226/GND (-2585 , 715.5)
*       104 = UAC116/U220/Gnd (-2577.5 , 667.5)
*       104 = UAC58/U238/B (-51.5 , 566.5)
*       104 = UAC58/U220/A (94 , 610.5)
*       104 = UAC58/U206/Gnd (131 , 595.5)
*       104 = UAC58/U220/GND (129 , 598)
*       104 = UAC58/U235/GND (183.5 , 554)
*       104 = UAC58/U229/Gnd (114 , 554.5)
*       104 = UAC90/U245/Gnd (-2585.5 , 554.5)
*       104 = UAC90/U218/Gnd (-2558.5 , 551.5)
*       104 = UAC90/U262/GND (-2587 , 598)
*       104 = UAC90/U222/Gnd (-2565 , 595.5)
*       104 = UAC105/U238/A (-2638.5 , 80)
*       104 = UAC105/U219/A (-2638 , 124)
*       104 = UAC105/B6 (-2638.5 , 51)
*       104 = UAC105/U235/A (-2412 , 80)
*       104 = UAC99/B6 (-2644.5 , 212.5)
*       104 = UAC99/U238/A (-2644.5 , 241.5)
*       104 = UAC99/U219/A (-2644 , 285.5)
*       104 = UAC99/U235/A (-2418 , 241.5)
*       104 = UAC94/U238/A (-2644 , 404)
*       104 = UAC94/B6 (-2644 , 375)
*       104 = UAC94/U235/A (-2417.5 , 404)
*       104 = UAC94/U219/A (-2643.5 , 448)
*       104 = UAC61/U238/B (-52 , 404)
*       104 = UAC61/U220/A (93.5 , 448)
*       104 = UAC61/C6 (93.5 , 480)
*       104 = UAC61/U235/GND (183 , 391.5)
*       104 = UAC61/U229/Gnd (113.5 , 392)
*       104 = UAC61/U253/GND (132 , 349)
*       104 = UAC61/U247/Gnd (157.5 , 348)
*       104 = UAC61/U246/Gnd (205.5 , 348)
*       104 = UAC59/U236/GND (-864 , 391.5)
*       104 = UAC59/U246/Gnd (-886 , 348)
*       104 = UAC94/U254/Gnd (-2522 , 348)
*       104 = UAC94/U245/Gnd (-2586 , 392)
*       104 = UAC94/U218/Gnd (-2559 , 389)
*       104 = UAC106/U238/A (-3005.5 , 80)
*       104 = UAC106/U219/A (-3005 , 124)
*       104 = UAC106/B6 (-3005.5 , 51)
*       104 = UAC106/U235/A (-2779 , 80)
*       104 = UAC100/B6 (-3011.5 , 212.5)
*       104 = UAC100/U238/A (-3011.5 , 241.5)
*       104 = UAC100/U219/A (-3011 , 285.5)
*       104 = UAC100/U235/A (-2785 , 241.5)
*       104 = UAC95/U238/A (-3011 , 404)
*       104 = UAC95/B6 (-3011 , 375)
*       104 = UAC65/U238/B (-52.5 , 241.5)
*       104 = UAC65/U220/A (93 , 285.5)
*       104 = UAC65/C6 (93 , 317.5)
*       104 = UAC99/U245/Gnd (-2586.5 , 229.5)
*       104 = UAC99/U218/Gnd (-2559.5 , 226.5)
*       104 = UAC99/U262/GND (-2588 , 273)
*       104 = UAC99/U222/Gnd (-2566 , 270.5)
*       104 = UAC107/U238/A (-3377 , 80)
*       104 = UAC107/U219/A (-3376.5 , 124)
*       104 = UAC107/B6 (-3377 , 51)
*       104 = UAC107/U235/A (-3150.5 , 80)
*       104 = UAC101/B6 (-3383 , 212.5)
*       104 = UAC70/U238/B (-53 , 80)
*       104 = UAC70/U220/A (92.5 , 124)
*       104 = UAC70/C6 (92.5 , 156)
*       104 = UAC62/U246/Gnd (-886.5 , 185.5)
*       104 = UAC68/U206/Gnd (-598.5 , 109)
*       104 = UAC68/U220/GND (-600.5 , 111.5)
*       104 = UAC68/U229/Gnd (-615.5 , 68)
*       104 = UAC68/U254/Gnd (-685.5 , 25.497)
*       104 = UAC109/U254/Gnd (-3627.5 , 24)
*       104 = UAC109/U253/GND (-3539 , 25)
*       104 = UAC109/U247/Gnd (-3513.5 , 24)
*       104 = UAC109/U246/Gnd (-3465.5 , 24)
*       104 = UAC107/U254/Gnd (-3255 , 24)
*       104 = UAC107/U253/GND (-3166.5 , 25)
*       104 = UAC107/U247/Gnd (-3141 , 24)
*       104 = UAC107/U246/Gnd (-3093 , 24)
*       104 = UAC106/U254/Gnd (-2883.5 , 24)
*       104 = UAC106/U253/GND (-2795 , 25)
*       104 = UAC106/U247/Gnd (-2769.5 , 24)
*       104 = UAC106/U246/Gnd (-2721.5 , 24)
*       104 = UAC105/U254/Gnd (-2516.5 , 24)
*       104 = UAC105/U253/GND (-2428 , 25)
*       104 = UAC105/U247/Gnd (-2402.5 , 24)
*       104 = UAC105/U246/Gnd (-2354.5 , 24)
*       104 = UAC104/U254/Gnd (-2146 , 24)
*       104 = UAC104/U253/GND (-2057.5 , 25)
*       104 = UAC104/U247/Gnd (-2032 , 24)
*       104 = UAC104/U246/Gnd (-1984 , 24)
*       104 = UAC103/U254/Gnd (-1782 , 24)
*       104 = UAC103/U253/GND (-1693.5 , 25)
*       104 = UAC103/U247/Gnd (-1668 , 24)
*       104 = UAC103/U246/Gnd (-1620 , 24)
*       104 = UAC102/U254/Gnd (-1414 , 24)
*       104 = UAC102/U253/GND (-1325.5 , 25)
*       104 = UAC102/U247/Gnd (-1300 , 24)
*       104 = UAC102/U246/Gnd (-1252 , 24)
*       104 = UAC67/U254/Gnd (-1049 , 24)
*       104 = UAC67/U253/GND (-960.5 , 25)
*       104 = UAC67/U247/Gnd (-935 , 24)
*       104 = UAC67/U246/Gnd (-887 , 24)
*       104 = UAC68/U253/GND (-597 , 25)
*       104 = UAC68/U247/Gnd (-571.5 , 24)
*       104 = UAC68/U246/Gnd (-523.5 , 24)
*       104 = UAC69/U254/Gnd (-321 , 24)
*       104 = UAC69/U253/GND (-232.5 , 25)
*       104 = UAC69/U247/Gnd (-207 , 24)
*       104 = UAC69/U246/Gnd (-159 , 24)
*       104 = UAC70/U254/Gnd (42.5 , 24)
*       104 = UAC70/U253/GND (131 , 25)
*       104 = UAC70/U247/Gnd (156.5 , 24)
*       104 = UAC70/U246/Gnd (204.5 , 24)
*       104 = UAC121/U230/GND (-3917.5 , 66.5)
*       104 = UAC121/U229/GND (-3934.5 , 66)
*       104 = UAC121/U228/GND (-3938.5 , 112)
*       104 = UAC121/U227/GND (-3964 , 112)
*       104 = UAC74/U238/B (-53.5 , -82.5)
*       104 = UAC74/U220/A (92 , -38.5)
*       104 = UAC74/C6 (92 , -6.5)
*       104 = UAC121/U220/Gnd (-3994 , 18.5)
*       104 = UAC121/U232/GND (-4022.5 , 21.5)
*       104 = UAC121/U231/GND (-4039.5 , 21)
*       104 = UAC73/U254/Gnd (-321.5 , -138.5)
*       104 = UAC73/U245/Gnd (-385.5 , -94.5)
*       104 = UAC73/U218/Gnd (-358.5 , -97.5)
*       104 = UAC72/U229/Gnd (-616 , -94.5)
*       104 = UAC72/U254/Gnd (-686 , -138.5)
*       104 = UAC72/U253/GND (-597.5 , -137.5)
*       104 = UAC71/U245/Gnd (-1113.5 , -94.5)
*       104 = UAC71/U238/GND (-1136.5 , -95)
*       104 = UAC71/U254/Gnd (-1049.5 , -138.5)
*       104 = UAC71/U218/Gnd (-1086.5 , -97.5)
*       104 = UAC71/U235/GND (-910 , -95)
*       104 = UAC71/U229/Gnd (-979.5 , -94.5)
*       104 = UAC71/U253/GND (-961 , -137.5)
*       104 = UAC71/U247/Gnd (-935.5 , -138.5)
*       104 = UAC71/U236/GND (-865.5 , -95)
*       104 = UAC71/U246/Gnd (-887.5 , -138.5)
*       104 = UAC72/U245/Gnd (-750 , -94.5)
*       104 = UAC72/U238/GND (-773 , -95)
*       104 = UAC72/U218/Gnd (-723 , -97.5)
*       104 = UAC72/U236/GND (-502 , -95)
*       104 = UAC72/U235/GND (-546.5 , -95)
*       104 = UAC72/U247/Gnd (-572 , -138.5)
*       104 = UAC72/U246/Gnd (-524 , -138.5)
*       104 = UAC73/U238/GND (-408.5 , -95)
*       104 = UAC73/U229/Gnd (-251.5 , -94.5)
*       104 = UAC73/U253/GND (-233 , -137.5)
*       104 = UAC73/U247/Gnd (-207.5 , -138.5)
*       104 = UAC73/U236/GND (-137.5 , -95)
*       104 = UAC73/U235/GND (-182 , -95)
*       104 = UAC73/U246/Gnd (-159.5 , -138.5)
*       104 = UAC74/U245/Gnd (-22 , -94.5)
*       104 = UAC74/U238/GND (-45 , -95)
*       104 = UAC74/U218/Gnd (5 , -97.5)
*       104 = UAC74/U254/Gnd (42 , -138.5)
*       104 = UAC74/U235/GND (181.5 , -95)
*       104 = UAC74/U229/Gnd (112 , -94.5)
*       104 = UAC74/U253/GND (130.5 , -137.5)
*       104 = UAC74/U247/Gnd (156 , -138.5)
*       104 = UAC74/U246/Gnd (204 , -138.5)
*       104 = UAC74/U236/GND (226 , -95)
*       104 = UAC126/Gnd (-1343 , -50.5)
*       104 = UAC125/GND (-1272 , -51)
*       104 = UAC124/Gnd (-1249 , -50.5)
*       104 = UAC71/F (-1209 , -30)
*       104 = UAC71/U262/GND (-1115 , -51)
*       104 = UAC71/U222/Gnd (-1093 , -53.5)
*       104 = UAC71/U219/GND (-1136 , -51)
*       104 = UAC71/U206/Gnd (-962.5 , -53.5)
*       104 = UAC71/U220/GND (-964.5 , -51)
*       104 = UAC72/F (-845.5 , -30)
*       104 = UAC71/U206/B (-885.5 , -38.5)
*       104 = UAC71/F6 (-881.5 , -10)
*       104 = UAC72/U262/GND (-751.5 , -51)
*       104 = UAC72/U222/Gnd (-729.5 , -53.5)
*       104 = UAC72/U219/GND (-772.5 , -51)
*       104 = UAC72/U206/Gnd (-599 , -53.5)
*       104 = UAC72/U220/GND (-601 , -51)
*       104 = UAC72/U206/B (-522 , -38.5)
*       104 = UAC72/F6 (-518 , -10)
*       104 = UAC73/U219/GND (-408 , -51)
*       104 = UAC73/F (-481 , -30)
*       104 = UAC73/U262/GND (-387 , -51)
*       104 = UAC73/U222/Gnd (-365 , -53.5)
*       104 = UAC73/U206/Gnd (-234.5 , -53.5)
*       104 = UAC73/U220/GND (-236.5 , -51)
*       104 = UAC74/F (-117.5 , -30)
*       104 = UAC73/U206/B (-157.5 , -38.5)
*       104 = UAC73/F6 (-153.5 , -10)
*       104 = UAC74/U262/GND (-23.5 , -51)
*       104 = UAC74/U222/Gnd (-1.5 , -53.5)
*       104 = UAC74/U219/GND (-44.5 , -51)
*       104 = UAC74/U206/Gnd (129 , -53.5)
*       104 = UAC74/U220/GND (127 , -51)
*       104 = UAC74/U206/B (206 , -38.5)
*       104 = UAC74/F6 (210 , -10)
*       104 = UAC74/U236/B (217.5 , -82.5)
*       104 = UAC74/C (258 , -55.5)
*       104 = UAC121/U223/GND (-4030.5 , 112)
*       104 = UAC121/U222/GND (-4047.5 , 111.5)
*       104 = UAC121/U226/GND (-4001.5 , 66.5)
*       104 = UAC121/U225/GND (-4018.5 , 66)
*       104 = UAC121/U224/GND (-4085.5 , 66.5)
*       104 = UAC109/U262/GND (-3693 , 111.5)
*       104 = UAC109/U245/Gnd (-3691.5 , 68)
*       104 = UAC109/U238/GND (-3714.5 , 67.5)
*       104 = UAC109/U219/GND (-3714 , 111.5)
*       104 = UAC109/U238/A (-3749.5 , 80)
*       104 = UAC109/U219/A (-3749 , 124)
*       104 = UAC109/B6 (-3749.5 , 51)
*       104 = UAC109/U218/Gnd (-3664.5 , 65)
*       104 = UAC109/U222/Gnd (-3671 , 109)
*       104 = UAC109/U206/Gnd (-3540.5 , 109)
*       104 = UAC109/U220/GND (-3542.5 , 111.5)
*       104 = UAC109/U229/Gnd (-3557.5 , 68)
*       104 = UAC109/U235/A (-3523 , 80)
*       104 = UAC109/U236/GND (-3443.5 , 67.5)
*       104 = UAC109/U235/GND (-3488 , 67.5)
*       104 = UAC107/U262/GND (-3320.5 , 111.5)
*       104 = UAC107/U222/Gnd (-3298.5 , 109)
*       104 = UAC107/U219/GND (-3341.5 , 111.5)
*       104 = UAC107/U245/Gnd (-3319 , 68)
*       104 = UAC107/U238/GND (-3342 , 67.5)
*       104 = UAC107/U218/Gnd (-3292 , 65)
*       104 = UAC107/U206/Gnd (-3168 , 109)
*       104 = UAC107/U220/GND (-3170 , 111.5)
*       104 = UAC107/U235/GND (-3115.5 , 67.5)
*       104 = UAC107/U229/Gnd (-3185 , 68)
*       104 = UAC107/U236/GND (-3071 , 67.5)
*       104 = UAC106/U245/Gnd (-2947.5 , 68)
*       104 = UAC106/U238/GND (-2970.5 , 67.5)
*       104 = UAC106/U218/Gnd (-2920.5 , 65)
*       104 = UAC106/U262/GND (-2949 , 111.5)
*       104 = UAC106/U222/Gnd (-2927 , 109)
*       104 = UAC106/U219/GND (-2970 , 111.5)
*       104 = UAC106/U206/Gnd (-2796.5 , 109)
*       104 = UAC106/U220/GND (-2798.5 , 111.5)
*       104 = UAC106/U229/Gnd (-2813.5 , 68)
*       104 = UAC106/U236/GND (-2699.5 , 67.5)
*       104 = UAC106/U235/GND (-2744 , 67.5)
*       104 = UAC105/U238/GND (-2603.5 , 67.5)
*       104 = UAC105/U219/GND (-2603 , 111.5)
*       104 = UAC105/U245/Gnd (-2580.5 , 68)
*       104 = UAC105/U218/Gnd (-2553.5 , 65)
*       104 = UAC105/U262/GND (-2582 , 111.5)
*       104 = UAC105/U222/Gnd (-2560 , 109)
*       104 = UAC105/U206/Gnd (-2429.5 , 109)
*       104 = UAC105/U220/GND (-2431.5 , 111.5)
*       104 = UAC105/U229/Gnd (-2446.5 , 68)
*       104 = UAC105/U236/GND (-2332.5 , 67.5)
*       104 = UAC105/U235/GND (-2377 , 67.5)
*       104 = UAC104/U262/GND (-2211.5 , 111.5)
*       104 = UAC104/U245/Gnd (-2210 , 68)
*       104 = UAC104/U238/GND (-2233 , 67.5)
*       104 = UAC104/U219/GND (-2232.5 , 111.5)
*       104 = UAC104/U218/Gnd (-2183 , 65)
*       104 = UAC104/U222/Gnd (-2189.5 , 109)
*       104 = UAC104/U206/Gnd (-2059 , 109)
*       104 = UAC104/U220/GND (-2061 , 111.5)
*       104 = UAC104/U235/GND (-2006.5 , 67.5)
*       104 = UAC104/U229/Gnd (-2076 , 68)
*       104 = UAC104/U236/GND (-1962 , 67.5)
*       104 = UAC103/U245/Gnd (-1846 , 68)
*       104 = UAC103/U238/GND (-1869 , 67.5)
*       104 = UAC103/U218/Gnd (-1819 , 65)
*       104 = UAC103/U262/GND (-1847.5 , 111.5)
*       104 = UAC103/U222/Gnd (-1825.5 , 109)
*       104 = UAC103/U219/GND (-1868.5 , 111.5)
*       104 = UAC103/U206/Gnd (-1695 , 109)
*       104 = UAC103/U220/GND (-1697 , 111.5)
*       104 = UAC103/U229/Gnd (-1712 , 68)
*       104 = UAC103/U236/GND (-1598 , 67.5)
*       104 = UAC103/U235/GND (-1642.5 , 67.5)
*       104 = UAC102/U238/GND (-1501 , 67.5)
*       104 = UAC102/U219/GND (-1500.5 , 111.5)
*       104 = UAC102/U245/Gnd (-1478 , 68)
*       104 = UAC102/U218/Gnd (-1451 , 65)
*       104 = UAC102/U262/GND (-1479.5 , 111.5)
*       104 = UAC102/U222/Gnd (-1457.5 , 109)
*       104 = UAC102/U206/Gnd (-1327 , 109)
*       104 = UAC102/U220/GND (-1329 , 111.5)
*       104 = UAC102/U229/Gnd (-1344 , 68)
*       104 = UAC102/U236/GND (-1230 , 67.5)
*       104 = UAC102/U235/GND (-1274.5 , 67.5)
*       104 = UAC67/U262/GND (-1114.5 , 111.5)
*       104 = UAC67/U222/Gnd (-1092.5 , 109)
*       104 = UAC67/U219/GND (-1135.5 , 111.5)
*       104 = UAC67/U245/Gnd (-1113 , 68)
*       104 = UAC67/U238/GND (-1136 , 67.5)
*       104 = UAC67/U218/Gnd (-1086 , 65)
*       104 = UAC67/U206/Gnd (-962 , 109)
*       104 = UAC67/U220/GND (-964 , 111.5)
*       104 = UAC67/U235/GND (-909.5 , 67.5)
*       104 = UAC67/U229/Gnd (-979 , 68)
*       104 = UAC67/U236/GND (-865 , 67.5)
*       104 = UAC68/U245/Gnd (-749.5 , 68)
*       104 = UAC68/U238/GND (-772.5 , 67.5)
*       104 = UAC68/U218/Gnd (-722.5 , 65)
*       104 = UAC68/U262/GND (-751 , 111.5)
*       104 = UAC68/U222/Gnd (-729 , 109)
*       104 = UAC68/U219/GND (-772 , 111.5)
*       104 = UAC68/U236/GND (-501.5 , 67.5)
*       104 = UAC68/U235/GND (-546 , 67.5)
*       104 = UAC69/U238/GND (-408 , 67.5)
*       104 = UAC69/U219/GND (-407.5 , 111.5)
*       104 = UAC69/U245/Gnd (-385 , 68)
*       104 = UAC69/U218/Gnd (-358 , 65)
*       104 = UAC69/U262/GND (-386.5 , 111.5)
*       104 = UAC69/U222/Gnd (-364.5 , 109)
*       104 = UAC69/U206/Gnd (-234 , 109)
*       104 = UAC69/U220/GND (-236 , 111.5)
*       104 = UAC69/U229/Gnd (-251 , 68)
*       104 = UAC69/U236/GND (-137 , 67.5)
*       104 = UAC69/U235/GND (-181.5 , 67.5)
*       104 = UAC70/U262/GND (-23 , 111.5)
*       104 = UAC70/U222/Gnd (-1 , 109)
*       104 = UAC70/U219/GND (-44 , 111.5)
*       104 = UAC70/U245/Gnd (-21.5 , 68)
*       104 = UAC70/U238/GND (-44.5 , 67.5)
*       104 = UAC70/U218/Gnd (5.5 , 65)
*       104 = UAC70/U206/Gnd (129.5 , 109)
*       104 = UAC70/U220/GND (127.5 , 111.5)
*       104 = UAC70/U235/GND (182 , 67.5)
*       104 = UAC70/U229/Gnd (112.5 , 68)
*       104 = UAC70/U236/GND (226.5 , 67.5)
*       104 = UAC70/U236/B (218 , 80)
*       104 = UAC70/C (258.5 , 107)
*       104 = UAC120/U232/GND (-3711.5 , 183)
*       104 = UAC120/U231/GND (-3728.5 , 182.5)
*       104 = UAC120/U220/Gnd (-3683 , 180)
*       104 = UAC101/U254/Gnd (-3261 , 185.5)
*       104 = UAC101/U253/GND (-3172.5 , 186.5)
*       104 = UAC101/U247/Gnd (-3147 , 185.5)
*       104 = UAC101/U246/Gnd (-3099 , 185.5)
*       104 = UAC100/U254/Gnd (-2889.5 , 185.5)
*       104 = UAC100/U253/GND (-2801 , 186.5)
*       104 = UAC100/U247/Gnd (-2775.5 , 185.5)
*       104 = UAC100/U246/Gnd (-2727.5 , 185.5)
*       104 = UAC99/U254/Gnd (-2522.5 , 185.5)
*       104 = UAC99/U253/GND (-2434 , 186.5)
*       104 = UAC99/U247/Gnd (-2408.5 , 185.5)
*       104 = UAC99/U246/Gnd (-2360.5 , 185.5)
*       104 = UAC98/U254/Gnd (-2152 , 185.5)
*       104 = UAC98/U253/GND (-2063.5 , 186.5)
*       104 = UAC98/U247/Gnd (-2038 , 185.5)
*       104 = UAC98/U246/Gnd (-1990 , 185.5)
*       104 = UAC97/U254/Gnd (-1788 , 185.5)
*       104 = UAC97/U253/GND (-1699.5 , 186.5)
*       104 = UAC97/U247/Gnd (-1674 , 185.5)
*       104 = UAC97/U246/Gnd (-1626 , 185.5)
*       104 = UAC96/U254/Gnd (-1420 , 185.5)
*       104 = UAC96/U253/GND (-1331.5 , 186.5)
*       104 = UAC96/U247/Gnd (-1306 , 185.5)
*       104 = UAC96/U246/Gnd (-1258 , 185.5)
*       104 = UAC62/U254/Gnd (-1048.5 , 185.5)
*       104 = UAC62/U253/GND (-960 , 186.5)
*       104 = UAC62/U247/Gnd (-934.5 , 185.5)
*       104 = UAC63/U254/Gnd (-685 , 185.5)
*       104 = UAC63/U253/GND (-596.5 , 186.5)
*       104 = UAC63/U247/Gnd (-571 , 185.5)
*       104 = UAC63/U246/Gnd (-523 , 185.5)
*       104 = UAC64/U254/Gnd (-320.5 , 185.5)
*       104 = UAC64/U253/GND (-232 , 186.5)
*       104 = UAC64/U247/Gnd (-206.5 , 185.5)
*       104 = UAC64/U246/Gnd (-158.5 , 185.5)
*       104 = UAC65/U254/Gnd (43 , 185.5)
*       104 = UAC65/U253/GND (131.5 , 186.5)
*       104 = UAC65/U247/Gnd (157 , 185.5)
*       104 = UAC65/U246/Gnd (205 , 185.5)
*       104 = UAC120/U223/GND (-3719.5 , 273.5)
*       104 = UAC120/U222/GND (-3736.5 , 273)
*       104 = UAC120/U225/GND (-3707.5 , 227.5)
*       104 = UAC120/U224/GND (-3774.5 , 228)
*       104 = UAC120/U230/GND (-3606.5 , 228)
*       104 = UAC120/U229/GND (-3623.5 , 227.5)
*       104 = UAC120/U226/GND (-3690.5 , 228)
*       104 = UAC120/U228/GND (-3627.5 , 273.5)
*       104 = UAC120/U227/GND (-3653 , 273.5)
*       104 = UAC101/U245/Gnd (-3325 , 229.5)
*       104 = UAC101/U238/GND (-3348 , 229)
*       104 = UAC101/U218/Gnd (-3298 , 226.5)
*       104 = UAC101/U262/GND (-3326.5 , 273)
*       104 = UAC101/U222/Gnd (-3304.5 , 270.5)
*       104 = UAC101/U219/GND (-3347.5 , 273)
*       104 = UAC101/U238/A (-3383 , 241.5)
*       104 = UAC101/U219/A (-3382.5 , 285.5)
*       104 = UAC101/U206/Gnd (-3174 , 270.5)
*       104 = UAC101/U220/GND (-3176 , 273)
*       104 = UAC101/U235/GND (-3121.5 , 229)
*       104 = UAC101/U229/Gnd (-3191 , 229.5)
*       104 = UAC101/U235/A (-3156.5 , 241.5)
*       104 = UAC101/U236/GND (-3077 , 229)
*       104 = UAC100/U245/Gnd (-2953.5 , 229.5)
*       104 = UAC100/U238/GND (-2976.5 , 229)
*       104 = UAC100/U218/Gnd (-2926.5 , 226.5)
*       104 = UAC100/U262/GND (-2955 , 273)
*       104 = UAC100/U222/Gnd (-2933 , 270.5)
*       104 = UAC100/U219/GND (-2976 , 273)
*       104 = UAC100/U206/Gnd (-2802.5 , 270.5)
*       104 = UAC100/U220/GND (-2804.5 , 273)
*       104 = UAC100/U229/Gnd (-2819.5 , 229.5)
*       104 = UAC100/U236/GND (-2705.5 , 229)
*       104 = UAC100/U235/GND (-2750 , 229)
*       104 = UAC99/U238/GND (-2609.5 , 229)
*       104 = UAC99/U219/GND (-2609 , 273)
*       104 = UAC99/U206/Gnd (-2435.5 , 270.5)
*       104 = UAC99/U220/GND (-2437.5 , 273)
*       104 = UAC99/U229/Gnd (-2452.5 , 229.5)
*       104 = UAC99/U236/GND (-2338.5 , 229)
*       104 = UAC99/U235/GND (-2383 , 229)
*       104 = UAC98/U262/GND (-2217.5 , 273)
*       104 = UAC98/U222/Gnd (-2195.5 , 270.5)
*       104 = UAC98/U219/GND (-2238.5 , 273)
*       104 = UAC98/U245/Gnd (-2216 , 229.5)
*       104 = UAC98/U238/GND (-2239 , 229)
*       104 = UAC98/U218/Gnd (-2189 , 226.5)
*       104 = UAC98/U206/Gnd (-2065 , 270.5)
*       104 = UAC98/U220/GND (-2067 , 273)
*       104 = UAC98/U235/GND (-2012.5 , 229)
*       104 = UAC98/U229/Gnd (-2082 , 229.5)
*       104 = UAC98/U236/GND (-1968 , 229)
*       104 = UAC97/U245/Gnd (-1852 , 229.5)
*       104 = UAC97/U238/GND (-1875 , 229)
*       104 = UAC97/U218/Gnd (-1825 , 226.5)
*       104 = UAC97/U262/GND (-1853.5 , 273)
*       104 = UAC97/U222/Gnd (-1831.5 , 270.5)
*       104 = UAC97/U219/GND (-1874.5 , 273)
*       104 = UAC97/U206/Gnd (-1701 , 270.5)
*       104 = UAC97/U220/GND (-1703 , 273)
*       104 = UAC97/U229/Gnd (-1718 , 229.5)
*       104 = UAC97/U236/GND (-1604 , 229)
*       104 = UAC97/U235/GND (-1648.5 , 229)
*       104 = UAC96/U238/GND (-1507 , 229)
*       104 = UAC96/U219/GND (-1506.5 , 273)
*       104 = UAC96/U245/Gnd (-1484 , 229.5)
*       104 = UAC96/U218/Gnd (-1457 , 226.5)
*       104 = UAC96/U262/GND (-1485.5 , 273)
*       104 = UAC96/U222/Gnd (-1463.5 , 270.5)
*       104 = UAC96/U206/Gnd (-1333 , 270.5)
*       104 = UAC96/U220/GND (-1335 , 273)
*       104 = UAC96/U229/Gnd (-1350 , 229.5)
*       104 = UAC96/U236/GND (-1236 , 229)
*       104 = UAC96/U235/GND (-1280.5 , 229)
*       104 = UAC62/U262/GND (-1114 , 273)
*       104 = UAC62/U245/Gnd (-1112.5 , 229.5)
*       104 = UAC62/U238/GND (-1135.5 , 229)
*       104 = UAC62/U222/Gnd (-1092 , 270.5)
*       104 = UAC62/U219/GND (-1135 , 273)
*       104 = UAC62/U218/Gnd (-1085.5 , 226.5)
*       104 = UAC62/U206/Gnd (-961.5 , 270.5)
*       104 = UAC62/U220/GND (-963.5 , 273)
*       104 = UAC62/U235/GND (-909 , 229)
*       104 = UAC62/U229/Gnd (-978.5 , 229.5)
*       104 = UAC62/U236/GND (-864.5 , 229)
*       104 = UAC63/U245/Gnd (-749 , 229.5)
*       104 = UAC63/U238/GND (-772 , 229)
*       104 = UAC63/U218/Gnd (-722 , 226.5)
*       104 = UAC63/U262/GND (-750.5 , 273)
*       104 = UAC63/U222/Gnd (-728.5 , 270.5)
*       104 = UAC63/U219/GND (-771.5 , 273)
*       104 = UAC63/U206/Gnd (-598 , 270.5)
*       104 = UAC63/U220/GND (-600 , 273)
*       104 = UAC63/U229/Gnd (-615 , 229.5)
*       104 = UAC63/U236/GND (-501 , 229)
*       104 = UAC63/U235/GND (-545.5 , 229)
*       104 = UAC64/U238/GND (-407.5 , 229)
*       104 = UAC64/U219/GND (-407 , 273)
*       104 = UAC64/U245/Gnd (-384.5 , 229.5)
*       104 = UAC64/U218/Gnd (-357.5 , 226.5)
*       104 = UAC64/U262/GND (-386 , 273)
*       104 = UAC64/U222/Gnd (-364 , 270.5)
*       104 = UAC64/U206/Gnd (-233.5 , 270.5)
*       104 = UAC64/U220/GND (-235.5 , 273)
*       104 = UAC64/U229/Gnd (-250.5 , 229.5)
*       104 = UAC64/U236/GND (-136.5 , 229)
*       104 = UAC64/U235/GND (-181 , 229)
*       104 = UAC65/U262/GND (-22.5 , 273)
*       104 = UAC65/U222/Gnd (-0.5 , 270.5)
*       104 = UAC65/U219/GND (-43.5 , 273)
*       104 = UAC65/U245/Gnd (-21 , 229.5)
*       104 = UAC65/U238/GND (-44 , 229)
*       104 = UAC65/U218/Gnd (6 , 226.5)
*       104 = UAC65/U206/Gnd (130 , 270.5)
*       104 = UAC65/U220/GND (128 , 273)
*       104 = UAC65/U235/GND (182.5 , 229)
*       104 = UAC65/U229/Gnd (113 , 229.5)
*       104 = UAC65/U236/GND (227 , 229)
*       104 = UAC65/U236/B (218.5 , 241.5)
*       104 = UAC65/C (259 , 268.5)
*       104 = UAC119/U224/GND (-3409.5 , 390.5)
*       104 = UAC119/U226/GND (-3325.5 , 390.5)
*       104 = UAC119/U225/GND (-3342.5 , 390)
*       104 = UAC119/U220/Gnd (-3318 , 342.5)
*       104 = UAC119/U232/GND (-3346.5 , 345.5)
*       104 = UAC119/U231/GND (-3363.5 , 345)
*       104 = UAC119/U230/GND (-3241.5 , 390.5)
*       104 = UAC119/U229/GND (-3258.5 , 390)
*       104 = UAC95/U245/Gnd (-2953 , 392)
*       104 = UAC95/U238/GND (-2976 , 391.5)
*       104 = UAC95/U218/Gnd (-2926 , 389)
*       104 = UAC95/U229/Gnd (-2819 , 392)
*       104 = UAC95/U254/Gnd (-2889 , 348)
*       104 = UAC95/U253/GND (-2800.5 , 349)
*       104 = UAC95/U236/GND (-2705 , 391.5)
*       104 = UAC95/U235/GND (-2749.5 , 391.5)
*       104 = UAC95/U247/Gnd (-2775 , 348)
*       104 = UAC95/U246/Gnd (-2727 , 348)
*       104 = UAC95/U235/A (-2784.5 , 404)
*       104 = UAC94/U238/GND (-2609 , 391.5)
*       104 = UAC94/U229/Gnd (-2452 , 392)
*       104 = UAC94/U253/GND (-2433.5 , 349)
*       104 = UAC94/U247/Gnd (-2408 , 348)
*       104 = UAC94/U236/GND (-2338 , 391.5)
*       104 = UAC94/U235/GND (-2382.5 , 391.5)
*       104 = UAC94/U246/Gnd (-2360 , 348)
*       104 = UAC93/U245/Gnd (-2215.5 , 392)
*       104 = UAC93/U238/GND (-2238.5 , 391.5)
*       104 = UAC93/U254/Gnd (-2151.5 , 348)
*       104 = UAC93/U218/Gnd (-2188.5 , 389)
*       104 = UAC93/U235/GND (-2012 , 391.5)
*       104 = UAC93/U229/Gnd (-2081.5 , 392)
*       104 = UAC93/U253/GND (-2063 , 349)
*       104 = UAC93/U247/Gnd (-2037.5 , 348)
*       104 = UAC93/U236/GND (-1967.5 , 391.5)
*       104 = UAC93/U246/Gnd (-1989.5 , 348)
*       104 = UAC92/U245/Gnd (-1851.5 , 392)
*       104 = UAC92/U238/GND (-1874.5 , 391.5)
*       104 = UAC92/U218/Gnd (-1824.5 , 389)
*       104 = UAC92/U229/Gnd (-1717.5 , 392)
*       104 = UAC92/U254/Gnd (-1787.5 , 348)
*       104 = UAC92/U253/GND (-1699 , 349)
*       104 = UAC92/U236/GND (-1603.5 , 391.5)
*       104 = UAC92/U235/GND (-1648 , 391.5)
*       104 = UAC92/U247/Gnd (-1673.5 , 348)
*       104 = UAC92/U246/Gnd (-1625.5 , 348)
*       104 = UAC91/U238/GND (-1506.5 , 391.5)
*       104 = UAC91/U254/Gnd (-1419.5 , 348)
*       104 = UAC91/U245/Gnd (-1483.5 , 392)
*       104 = UAC91/U218/Gnd (-1456.5 , 389)
*       104 = UAC91/U229/Gnd (-1349.5 , 392)
*       104 = UAC91/U253/GND (-1331 , 349)
*       104 = UAC91/U247/Gnd (-1305.5 , 348)
*       104 = UAC91/U236/GND (-1235.5 , 391.5)
*       104 = UAC91/U235/GND (-1280 , 391.5)
*       104 = UAC91/U246/Gnd (-1257.5 , 348)
*       104 = UAC59/U245/Gnd (-1112 , 392)
*       104 = UAC59/U238/GND (-1135 , 391.5)
*       104 = UAC59/U254/Gnd (-1048 , 348)
*       104 = UAC59/U218/Gnd (-1085 , 389)
*       104 = UAC59/U235/GND (-908.5 , 391.5)
*       104 = UAC59/U229/Gnd (-978 , 392)
*       104 = UAC59/U253/GND (-959.5 , 349)
*       104 = UAC59/U247/Gnd (-934 , 348)
*       104 = UAC66/U245/Gnd (-748.5 , 392)
*       104 = UAC66/U238/GND (-771.5 , 391.5)
*       104 = UAC66/U218/Gnd (-721.5 , 389)
*       104 = UAC66/U229/Gnd (-614.5 , 392)
*       104 = UAC66/U254/Gnd (-684.5 , 348)
*       104 = UAC66/U253/GND (-596 , 349)
*       104 = UAC66/U236/GND (-500.5 , 391.5)
*       104 = UAC66/U235/GND (-545 , 391.5)
*       104 = UAC66/U247/Gnd (-570.5 , 348)
*       104 = UAC66/U246/Gnd (-522.5 , 348)
*       104 = UAC60/U238/GND (-407 , 391.5)
*       104 = UAC60/U254/Gnd (-320 , 348)
*       104 = UAC60/U245/Gnd (-384 , 392)
*       104 = UAC60/U218/Gnd (-357 , 389)
*       104 = UAC60/U229/Gnd (-250 , 392)
*       104 = UAC60/U253/GND (-231.5 , 349)
*       104 = UAC60/U247/Gnd (-206 , 348)
*       104 = UAC60/U236/GND (-136 , 391.5)
*       104 = UAC60/U235/GND (-180.5 , 391.5)
*       104 = UAC60/U246/Gnd (-158 , 348)
*       104 = UAC61/U245/Gnd (-20.5 , 392)
*       104 = UAC61/U238/GND (-43.5 , 391.5)
*       104 = UAC61/U218/Gnd (6.5 , 389)
*       104 = UAC61/U254/Gnd (43.5 , 348)
*       104 = UAC61/U236/GND (227.5 , 391.5)
*       104 = UAC119/U223/GND (-3354.5 , 436)
*       104 = UAC119/U222/GND (-3371.5 , 435.5)
*       104 = UAC119/U228/GND (-3262.5 , 436)
*       104 = UAC119/U227/GND (-3288 , 436)
*       104 = UAC95/U219/A (-3010.5 , 448)
*       104 = UAC95/U262/GND (-2954.5 , 435.5)
*       104 = UAC95/U222/Gnd (-2932.5 , 433)
*       104 = UAC95/U219/GND (-2975.5 , 435.5)
*       104 = UAC118/U220/Gnd (-2943.5 , 505)
*       104 = UAC118/U232/GND (-2972 , 508)
*       104 = UAC118/U231/GND (-2989 , 507.5)
*       104 = UAC95/U206/Gnd (-2802 , 433)
*       104 = UAC95/U220/GND (-2804 , 435.5)
*       104 = UAC94/U219/GND (-2608.5 , 435.5)
*       104 = UAC90/U254/Gnd (-2521.5 , 510.5)
*       104 = UAC94/U262/GND (-2587.5 , 435.5)
*       104 = UAC94/U222/Gnd (-2565.5 , 433)
*       104 = UAC90/U253/GND (-2433 , 511.5)
*       104 = UAC90/U247/Gnd (-2407.5 , 510.5)
*       104 = UAC94/U206/Gnd (-2435 , 433)
*       104 = UAC94/U220/GND (-2437 , 435.5)
*       104 = UAC90/U246/Gnd (-2359.5 , 510.5)
*       104 = UAC93/U262/GND (-2217 , 435.5)
*       104 = UAC93/U222/Gnd (-2195 , 433)
*       104 = UAC93/U219/GND (-2238 , 435.5)
*       104 = UAC88/U254/Gnd (-2151 , 510.5)
*       104 = UAC88/U253/GND (-2062.5 , 511.5)
*       104 = UAC88/U247/Gnd (-2037 , 510.5)
*       104 = UAC93/U206/Gnd (-2064.5 , 433)
*       104 = UAC93/U220/GND (-2066.5 , 435.5)
*       104 = UAC88/U246/Gnd (-1989 , 510.5)
*       104 = UAC92/U262/GND (-1853 , 435.5)
*       104 = UAC92/U222/Gnd (-1831 , 433)
*       104 = UAC92/U219/GND (-1874 , 435.5)
*       104 = UAC87/U254/Gnd (-1787 , 510.5)
*       104 = UAC87/U253/GND (-1698.5 , 511.5)
*       104 = UAC92/U206/Gnd (-1700.5 , 433)
*       104 = UAC92/U220/GND (-1702.5 , 435.5)
*       104 = UAC87/U247/Gnd (-1673 , 510.5)
*       104 = UAC87/U246/Gnd (-1625 , 510.5)
*       104 = UAC91/U219/GND (-1506 , 435.5)
*       104 = UAC85/U254/Gnd (-1419 , 510.5)
*       104 = UAC91/U262/GND (-1485 , 435.5)
*       104 = UAC91/U222/Gnd (-1463 , 433)
*       104 = UAC85/U253/GND (-1330.5 , 511.5)
*       104 = UAC85/U247/Gnd (-1305 , 510.5)
*       104 = UAC91/U206/Gnd (-1332.5 , 433)
*       104 = UAC91/U220/GND (-1334.5 , 435.5)
*       104 = UAC85/U246/Gnd (-1257 , 510.5)
*       104 = UAC59/U262/GND (-1113.5 , 435.5)
*       104 = UAC59/U222/Gnd (-1091.5 , 433)
*       104 = UAC59/U219/GND (-1134.5 , 435.5)
*       104 = UAC55/U254/Gnd (-1047.5 , 510.5)
*       104 = UAC55/U253/GND (-959 , 511.5)
*       104 = UAC55/U247/Gnd (-933.5 , 510.5)
*       104 = UAC59/U206/Gnd (-961 , 433)
*       104 = UAC59/U220/GND (-963 , 435.5)
*       104 = UAC55/U246/Gnd (-885.5 , 510.5)
*       104 = UAC66/U262/GND (-750 , 435.5)
*       104 = UAC66/U222/Gnd (-728 , 433)
*       104 = UAC66/U219/GND (-771 , 435.5)
*       104 = UAC56/U254/Gnd (-684 , 510.5)
*       104 = UAC56/U253/GND (-595.5 , 511.5)
*       104 = UAC66/U206/Gnd (-597.5 , 433)
*       104 = UAC66/U220/GND (-599.5 , 435.5)
*       104 = UAC56/U247/Gnd (-570 , 510.5)
*       104 = UAC56/U246/Gnd (-522 , 510.5)
*       104 = UAC60/U219/GND (-406.5 , 435.5)
*       104 = UAC57/U254/Gnd (-319.5 , 510.5)
*       104 = UAC60/U262/GND (-385.5 , 435.5)
*       104 = UAC60/U222/Gnd (-363.5 , 433)
*       104 = UAC57/U253/GND (-231 , 511.5)
*       104 = UAC57/U247/Gnd (-205.5 , 510.5)
*       104 = UAC60/U206/Gnd (-233 , 433)
*       104 = UAC60/U220/GND (-235 , 435.5)
*       104 = UAC57/U246/Gnd (-157.5 , 510.5)
*       104 = UAC61/U262/GND (-22 , 435.5)
*       104 = UAC61/U222/Gnd (0 , 433)
*       104 = UAC61/U219/GND (-43 , 435.5)
*       104 = UAC58/U254/Gnd (44 , 510.5)
*       104 = UAC58/U253/GND (132.5 , 511.5)
*       104 = UAC58/U247/Gnd (158 , 510.5)
*       104 = UAC58/U246/Gnd (206 , 510.5)
*       104 = UAC61/U206/Gnd (130.5 , 433)
*       104 = UAC61/U220/GND (128.5 , 435.5)
*       104 = UAC61/U236/B (219 , 404)
*       104 = UAC61/C (259.5 , 431)
*       104 = UAC118/U222/GND (-2997 , 598)
*       104 = UAC118/U224/GND (-3035 , 553)
*       104 = UAC118/U227/GND (-2913.5 , 598.5)
*       104 = UAC118/U223/GND (-2980 , 598.5)
*       104 = UAC118/U226/GND (-2951 , 553)
*       104 = UAC118/U225/GND (-2968 , 552.5)
*       104 = UAC118/U230/GND (-2867 , 553)
*       104 = UAC118/U229/GND (-2884 , 552.5)
*       104 = UAC118/U228/GND (-2888 , 598.5)
*       104 = UAC90/U238/GND (-2608.5 , 554)
*       104 = UAC90/U219/GND (-2608 , 598)
*       104 = UAC90/U238/A (-2643.5 , 566.5)
*       104 = UAC90/U219/A (-2643 , 610.5)
*       104 = UAC90/B6 (-2643.5 , 537.5)
*       104 = UAC90/U206/Gnd (-2434.5 , 595.5)
*       104 = UAC90/U220/GND (-2436.5 , 598)
*       104 = UAC90/U229/Gnd (-2451.5 , 554.5)
*       104 = UAC90/U235/A (-2417 , 566.5)
*       104 = UAC90/U236/GND (-2337.5 , 554)
*       104 = UAC90/U235/GND (-2382 , 554)
*       104 = UAC88/U262/GND (-2216.5 , 598)
*       104 = UAC88/U222/Gnd (-2194.5 , 595.5)
*       104 = UAC88/U219/GND (-2237.5 , 598)
*       104 = UAC88/U245/Gnd (-2215 , 554.5)
*       104 = UAC88/U238/GND (-2238 , 554)
*       104 = UAC88/U218/Gnd (-2188 , 551.5)
*       104 = UAC88/U206/Gnd (-2064 , 595.5)
*       104 = UAC88/U220/GND (-2066 , 598)
*       104 = UAC88/U235/GND (-2011.5 , 554)
*       104 = UAC88/U229/Gnd (-2081 , 554.5)
*       104 = UAC88/U236/GND (-1967 , 554)
*       104 = UAC87/U245/Gnd (-1851 , 554.5)
*       104 = UAC87/U238/GND (-1874 , 554)
*       104 = UAC87/U218/Gnd (-1824 , 551.5)
*       104 = UAC87/U262/GND (-1852.5 , 598)
*       104 = UAC87/U222/Gnd (-1830.5 , 595.5)
*       104 = UAC87/U219/GND (-1873.5 , 598)
*       104 = UAC87/U206/Gnd (-1700 , 595.5)
*       104 = UAC87/U220/GND (-1702 , 598)
*       104 = UAC87/U229/Gnd (-1717 , 554.5)
*       104 = UAC87/U236/GND (-1603 , 554)
*       104 = UAC87/U235/GND (-1647.5 , 554)
*       104 = UAC85/U238/GND (-1506 , 554)
*       104 = UAC85/U219/GND (-1505.5 , 598)
*       104 = UAC85/U245/Gnd (-1483 , 554.5)
*       104 = UAC85/U218/Gnd (-1456 , 551.5)
*       104 = UAC85/U262/GND (-1484.5 , 598)
*       104 = UAC85/U222/Gnd (-1462.5 , 595.5)
*       104 = UAC85/U206/Gnd (-1332 , 595.5)
*       104 = UAC85/U220/GND (-1334 , 598)
*       104 = UAC85/U229/Gnd (-1349 , 554.5)
*       104 = UAC85/U236/GND (-1235 , 554)
*       104 = UAC85/U235/GND (-1279.5 , 554)
*       104 = UAC55/U262/GND (-1113 , 598)
*       104 = UAC55/U245/Gnd (-1111.5 , 554.5)
*       104 = UAC55/U238/GND (-1134.5 , 554)
*       104 = UAC55/U219/GND (-1134 , 598)
*       104 = UAC55/U218/Gnd (-1084.5 , 551.5)
*       104 = UAC55/U222/Gnd (-1091 , 595.5)
*       104 = UAC55/U206/Gnd (-960.5 , 595.5)
*       104 = UAC55/U220/GND (-962.5 , 598)
*       104 = UAC55/U235/GND (-908 , 554)
*       104 = UAC55/U229/Gnd (-977.5 , 554.5)
*       104 = UAC55/U236/GND (-863.5 , 554)
*       104 = UAC56/U245/Gnd (-748 , 554.5)
*       104 = UAC56/U238/GND (-771 , 554)
*       104 = UAC56/U218/Gnd (-721 , 551.5)
*       104 = UAC56/U262/GND (-749.5 , 598)
*       104 = UAC56/U222/Gnd (-727.5 , 595.5)
*       104 = UAC56/U219/GND (-770.5 , 598)
*       104 = UAC56/U206/Gnd (-597 , 595.5)
*       104 = UAC56/U220/GND (-599 , 598)
*       104 = UAC56/U229/Gnd (-614 , 554.5)
*       104 = UAC56/U236/GND (-500 , 554)
*       104 = UAC56/U235/GND (-544.5 , 554)
*       104 = UAC57/U238/GND (-406.5 , 554)
*       104 = UAC57/U219/GND (-406 , 598)
*       104 = UAC57/U245/Gnd (-383.5 , 554.5)
*       104 = UAC57/U218/Gnd (-356.5 , 551.5)
*       104 = UAC57/U262/GND (-385 , 598)
*       104 = UAC57/U222/Gnd (-363 , 595.5)
*       104 = UAC57/U206/Gnd (-232.5 , 595.5)
*       104 = UAC57/U220/GND (-234.5 , 598)
*       104 = UAC57/U229/Gnd (-249.5 , 554.5)
*       104 = UAC57/U236/GND (-135.5 , 554)
*       104 = UAC57/U235/GND (-180 , 554)
*       104 = UAC58/U262/GND (-21.5 , 598)
*       104 = UAC58/U222/Gnd (0.5 , 595.5)
*       104 = UAC58/U219/GND (-42.5 , 598)
*       104 = UAC58/U245/Gnd (-20 , 554.5)
*       104 = UAC58/U238/GND (-43 , 554)
*       104 = UAC58/U218/Gnd (7 , 551.5)
*       104 = UAC58/U236/GND (228 , 554)
*       104 = UAC58/U236/B (219.5 , 566.5)
*       104 = UAC58/C (260 , 593.5)
*       104 = UAC116/U225/GND (-2602 , 715)
*       104 = UAC116/U224/GND (-2669 , 715.5)
*       104 = UAC116/U232/GND (-2606 , 670.5)
*       104 = UAC116/U231/GND (-2623 , 670)
*       104 = UAC84/U245/Gnd (-2214.5 , 717)
*       104 = UAC84/U238/GND (-2237.5 , 716.5)
*       104 = UAC84/B6 (-2272.5 , 700)
*       104 = UAC84/U254/Gnd (-2150.5 , 673)
*       104 = UAC84/U218/Gnd (-2187.5 , 714)
*       104 = UAC84/U235/GND (-2011 , 716.5)
*       104 = UAC84/U229/Gnd (-2080.5 , 717)
*       104 = UAC84/U253/GND (-2062 , 674)
*       104 = UAC84/U247/Gnd (-2036.5 , 673)
*       104 = UAC84/U236/GND (-1966.5 , 716.5)
*       104 = UAC84/U246/Gnd (-1988.5 , 673)
*       104 = UAC82/U245/Gnd (-1851 , 717)
*       104 = UAC82/U238/GND (-1874 , 716.5)
*       104 = UAC82/U218/Gnd (-1824 , 714)
*       104 = UAC82/U229/Gnd (-1717 , 717)
*       104 = UAC82/U254/Gnd (-1787 , 673)
*       104 = UAC82/U253/GND (-1698.5 , 674)
*       104 = UAC82/U236/GND (-1603 , 716.5)
*       104 = UAC82/U235/GND (-1647.5 , 716.5)
*       104 = UAC82/U247/Gnd (-1673 , 673)
*       104 = UAC82/U246/Gnd (-1625 , 673)
*       104 = UAC81/U238/GND (-1505.5 , 716.5)
*       104 = UAC81/U254/Gnd (-1418.5 , 673)
*       104 = UAC81/U245/Gnd (-1482.5 , 717)
*       104 = UAC81/U218/Gnd (-1455.5 , 714)
*       104 = UAC81/U229/Gnd (-1348.5 , 717)
*       104 = UAC81/U253/GND (-1330 , 674)
*       104 = UAC81/U247/Gnd (-1304.5 , 673)
*       104 = UAC81/U236/GND (-1234.5 , 716.5)
*       104 = UAC81/U235/GND (-1279 , 716.5)
*       104 = UAC81/U246/Gnd (-1256.5 , 673)
*       104 = UAC51/U245/Gnd (-1111 , 717)
*       104 = UAC51/U238/GND (-1134 , 716.5)
*       104 = UAC51/U254/Gnd (-1047 , 673)
*       104 = UAC51/U218/Gnd (-1084 , 714)
*       104 = UAC51/U235/GND (-907.5 , 716.5)
*       104 = UAC51/U229/Gnd (-977 , 717)
*       104 = UAC51/U253/GND (-958.5 , 674)
*       104 = UAC51/U247/Gnd (-933 , 673)
*       104 = UAC51/U236/GND (-863 , 716.5)
*       104 = UAC51/U246/Gnd (-885 , 673)
*       104 = UAC52/U245/Gnd (-747.5 , 717)
*       104 = UAC52/U238/GND (-770.5 , 716.5)
*       104 = UAC52/U218/Gnd (-720.5 , 714)
*       104 = UAC52/U229/Gnd (-613.5 , 717)
*       104 = UAC52/U254/Gnd (-683.5 , 673)
*       104 = UAC52/U253/GND (-595 , 674)
*       104 = UAC52/U236/GND (-499.5 , 716.5)
*       104 = UAC52/U235/GND (-544 , 716.5)
*       104 = UAC52/U247/Gnd (-569.5 , 673)
*       104 = UAC52/U246/Gnd (-521.5 , 673)
*       104 = UAC53/U238/GND (-406 , 716.5)
*       104 = UAC53/U254/Gnd (-319 , 673)
*       104 = UAC53/U245/Gnd (-383 , 717)
*       104 = UAC53/U218/Gnd (-356 , 714)
*       104 = UAC53/U229/Gnd (-249 , 717)
*       104 = UAC53/U253/GND (-230.5 , 674)
*       104 = UAC53/U247/Gnd (-205 , 673)
*       104 = UAC53/U236/GND (-135 , 716.5)
*       104 = UAC53/U235/GND (-179.5 , 716.5)
*       104 = UAC53/U246/Gnd (-157 , 673)
*       104 = UAC54/U245/Gnd (-19.5 , 717)
*       104 = UAC54/U238/GND (-42.5 , 716.5)
*       104 = UAC54/U218/Gnd (7.5 , 714)
*       104 = UAC54/U254/Gnd (44.5 , 673)
*       104 = UAC58/C6 (94 , 642.5)
*       104 = UAC54/U236/GND (228.5 , 716.5)
*       104 = UAC116/U223/GND (-2614 , 761)
*       104 = UAC116/U222/GND (-2631 , 760.5)
*       104 = UAC116/U228/GND (-2522 , 761)
*       104 = UAC116/U227/GND (-2547.5 , 761)
*       104 = UAC84/U262/GND (-2216 , 760.5)
*       104 = UAC84/U222/Gnd (-2194 , 758)
*       104 = UAC84/U219/GND (-2237 , 760.5)
*       104 = UAC84/U238/A (-2272.5 , 729)
*       104 = UAC84/U219/A (-2272 , 773)
*       104 = UAC84/U206/Gnd (-2063.5 , 758)
*       104 = UAC84/U220/GND (-2065.5 , 760.5)
*       104 = UAC84/U235/A (-2046 , 729)
*       104 = UAC82/U262/GND (-1852.5 , 760.5)
*       104 = UAC82/U222/Gnd (-1830.5 , 758)
*       104 = UAC82/U219/GND (-1873.5 , 760.5)
*       104 = UAC82/U206/Gnd (-1700 , 758)
*       104 = UAC82/U220/GND (-1702 , 760.5)
*       104 = UAC81/U219/GND (-1505 , 760.5)
*       104 = UAC81/U262/GND (-1484 , 760.5)
*       104 = UAC81/U222/Gnd (-1462 , 758)
*       104 = UAC81/U206/Gnd (-1331.5 , 758)
*       104 = UAC81/U220/GND (-1333.5 , 760.5)
*       104 = UAC51/U262/GND (-1112.5 , 760.5)
*       104 = UAC51/U219/GND (-1133.5 , 760.5)
*       104 = UAC51/U222/Gnd (-1090.5 , 758)
*       104 = UAC51/U206/Gnd (-960 , 758)
*       104 = UAC51/U220/GND (-962 , 760.5)
*       104 = UAC52/U262/GND (-749 , 760.5)
*       104 = UAC52/U222/Gnd (-727 , 758)
*       104 = UAC52/U219/GND (-770 , 760.5)
*       104 = UAC52/U206/Gnd (-596.5 , 758)
*       104 = UAC52/U220/GND (-598.5 , 760.5)
*       104 = UAC53/U219/GND (-405.5 , 760.5)
*       104 = UAC53/U262/GND (-384.5 , 760.5)
*       104 = UAC53/U222/Gnd (-362.5 , 758)
*       104 = UAC53/U206/Gnd (-232 , 758)
*       104 = UAC53/U220/GND (-234 , 760.5)
*       104 = UAC54/U262/GND (-21 , 760.5)
*       104 = UAC54/U222/Gnd (1 , 758)
*       104 = UAC54/U219/GND (-42 , 760.5)
*       104 = UAC54/U206/Gnd (131.5 , 758)
*       104 = UAC54/U220/GND (129.5 , 760.5)
*       104 = UAC54/U236/B (220 , 729)
*       104 = UAC54/C (260.5 , 756)
*       104 = UAC114/U226/GND (-2214 , 877)
*       104 = UAC114/U225/GND (-2231 , 876.5)
*       104 = UAC114/U220/Gnd (-2206.5 , 829)
*       104 = UAC114/U232/GND (-2235 , 832)
*       104 = UAC114/U231/GND (-2252 , 831.5)
*       104 = UAC114/U230/GND (-2130 , 877)
*       104 = UAC114/U229/GND (-2147 , 876.5)
*       104 = UAC114/U228/GND (-2151 , 922.5)
*       104 = UAC114/U227/GND (-2176.5 , 922.5)
*       104 = UAC103/U238/A (-1904 , 80)
*       104 = UAC103/U219/A (-1903.5 , 124)
*       104 = UAC103/B6 (-1904 , 51)
*       104 = UAC103/U235/A (-1677.5 , 80)
*       104 = UAC97/B6 (-1910 , 212.5)
*       104 = UAC97/U238/A (-1910 , 241.5)
*       104 = UAC97/U219/A (-1909.5 , 285.5)
*       104 = UAC97/U235/A (-1683.5 , 241.5)
*       104 = UAC92/U238/A (-1909.5 , 404)
*       104 = UAC92/B6 (-1909.5 , 375)
*       104 = UAC92/U235/A (-1683 , 404)
*       104 = UAC92/U219/A (-1909 , 448)
*       104 = UAC87/U238/A (-1909 , 566.5)
*       104 = UAC87/U219/A (-1908.5 , 610.5)
*       104 = UAC87/B6 (-1909 , 537.5)
*       104 = UAC87/U235/A (-1682.5 , 566.5)
*       104 = UAC82/B6 (-1909 , 700)
*       104 = UAC82/U238/A (-1909 , 729)
*       104 = UAC82/U219/A (-1908.5 , 773)
*       104 = UAC82/U235/A (-1682.5 , 729)
*       104 = UAC80/U238/A (-1896 , 890.5)
*       104 = UAC80/B6 (-1896 , 861.5)
*       104 = UAC80/U262/GND (-1839.5 , 922)
*       104 = UAC80/U222/Gnd (-1817.5 , 919.5)
*       104 = UAC80/U219/GND (-1860.5 , 922)
*       104 = UAC80/U245/Gnd (-1838 , 878.5)
*       104 = UAC80/U238/GND (-1861 , 878)
*       104 = UAC80/U218/Gnd (-1811 , 875.5)
*       104 = UAC80/U229/Gnd (-1704 , 878.5)
*       104 = UAC80/U254/Gnd (-1774 , 834.5)
*       104 = UAC80/U206/Gnd (-1687 , 919.5)
*       104 = UAC80/U220/GND (-1689 , 922)
*       104 = UAC80/U235/GND (-1634.5 , 878)
*       104 = UAC80/U253/GND (-1685.5 , 835.5)
*       104 = UAC80/U247/Gnd (-1660 , 834.5)
*       104 = UAC80/U246/Gnd (-1612 , 834.5)
*       104 = UAC80/U235/A (-1669.5 , 890.5)
*       104 = UAC80/U236/GND (-1590 , 878)
*       104 = UAC79/U238/GND (-1497.5 , 878)
*       104 = UAC79/U219/GND (-1497 , 922)
*       104 = UAC79/U262/GND (-1476 , 922)
*       104 = UAC79/U222/Gnd (-1454 , 919.5)
*       104 = UAC79/U254/Gnd (-1410.5 , 834.5)
*       104 = UAC79/U245/Gnd (-1474.5 , 878.5)
*       104 = UAC79/U218/Gnd (-1447.5 , 875.5)
*       104 = UAC79/U206/Gnd (-1323.5 , 919.5)
*       104 = UAC79/U220/GND (-1325.5 , 922)
*       104 = UAC79/U229/Gnd (-1340.5 , 878.5)
*       104 = UAC79/U253/GND (-1322 , 835.5)
*       104 = UAC79/U247/Gnd (-1296.5 , 834.5)
*       104 = UAC79/U236/GND (-1226.5 , 878)
*       104 = UAC79/U235/GND (-1271 , 878)
*       104 = UAC79/U246/Gnd (-1248.5 , 834.5)
*       104 = UAC39/U262/GND (-1112 , 922)
*       104 = UAC39/U245/Gnd (-1110.5 , 878.5)
*       104 = UAC39/U238/GND (-1133.5 , 878)
*       104 = UAC39/U219/GND (-1133 , 922)
*       104 = UAC39/U254/Gnd (-1046.5 , 834.5)
*       104 = UAC39/U218/Gnd (-1083.5 , 875.5)
*       104 = UAC39/U222/Gnd (-1090 , 919.5)
*       104 = UAC39/U206/Gnd (-959.5 , 919.5)
*       104 = UAC39/U220/GND (-961.5 , 922)
*       104 = UAC39/U235/GND (-907 , 878)
*       104 = UAC39/U229/Gnd (-976.5 , 878.5)
*       104 = UAC39/U253/GND (-958 , 835.5)
*       104 = UAC39/U247/Gnd (-932.5 , 834.5)
*       104 = UAC39/U236/GND (-862.5 , 878)
*       104 = UAC39/U246/Gnd (-884.5 , 834.5)
*       104 = UAC40/U245/Gnd (-747 , 878.5)
*       104 = UAC40/U238/GND (-770 , 878)
*       104 = UAC40/U218/Gnd (-720 , 875.5)
*       104 = UAC40/U206/Gnd (-596 , 919.5)
*       104 = UAC40/U220/GND (-598 , 922)
*       104 = UAC40/U229/Gnd (-613 , 878.5)
*       104 = UAC40/U254/Gnd (-683 , 834.5)
*       104 = UAC40/U253/GND (-594.5 , 835.5)
*       104 = UAC40/U236/GND (-499 , 878)
*       104 = UAC40/U235/GND (-543.5 , 878)
*       104 = UAC40/U247/Gnd (-569 , 834.5)
*       104 = UAC40/U246/Gnd (-521 , 834.5)
*       104 = UAC41/U238/GND (-405.5 , 878)
*       104 = UAC41/U219/GND (-405 , 922)
*       104 = UAC41/U262/GND (-384 , 922)
*       104 = UAC41/U222/Gnd (-362 , 919.5)
*       104 = UAC41/U254/Gnd (-318.5 , 834.5)
*       104 = UAC41/U245/Gnd (-382.5 , 878.5)
*       104 = UAC41/U218/Gnd (-355.5 , 875.5)
*       104 = UAC41/U206/Gnd (-231.5 , 919.5)
*       104 = UAC41/U220/GND (-233.5 , 922)
*       104 = UAC41/U229/Gnd (-248.5 , 878.5)
*       104 = UAC41/U253/GND (-230 , 835.5)
*       104 = UAC41/U247/Gnd (-204.5 , 834.5)
*       104 = UAC41/U236/GND (-134.5 , 878)
*       104 = UAC41/U235/GND (-179 , 878)
*       104 = UAC41/U246/Gnd (-156.5 , 834.5)
*       104 = UAC42/U245/Gnd (-19 , 878.5)
*       104 = UAC42/U238/GND (-42 , 878)
*       104 = UAC42/U218/Gnd (8 , 875.5)
*       104 = UAC42/U254/Gnd (45 , 834.5)
*       104 = UAC42/U206/Gnd (132 , 919.5)
*       104 = UAC42/U220/GND (130 , 922)
*       104 = UAC42/U235/GND (184.5 , 878)
*       104 = UAC42/U229/Gnd (115 , 878.5)
*       104 = UAC42/U253/GND (133.5 , 835.5)
*       104 = UAC42/U247/Gnd (159 , 834.5)
*       104 = UAC42/U246/Gnd (207 , 834.5)
*       104 = UAC42/U236/GND (229 , 878)
*       104 = UAC42/U236/B (220.5 , 890.5)
*       104 = UAC42/C (261 , 917.5)
*       104 = UAC80/U219/A (-1895.5 , 934.5)
*       104 = UAC112/U220/Gnd (-1829.5 , 991.5)
*       104 = UAC112/U232/GND (-1858 , 994.5)
*       104 = UAC112/U231/GND (-1875 , 994)
*       104 = UAC78/U254/Gnd (-1410 , 997)
*       104 = UAC78/U253/GND (-1321.5 , 998)
*       104 = UAC78/U247/Gnd (-1296 , 997)
*       104 = UAC78/U246/Gnd (-1248 , 997)
*       104 = UAC35/U254/Gnd (-1046 , 997)
*       104 = UAC35/U253/GND (-957.5 , 998)
*       104 = UAC35/U247/Gnd (-932 , 997)
*       104 = UAC35/U246/Gnd (-884 , 997)
*       104 = UAC36/U254/Gnd (-682.5 , 997)
*       104 = UAC36/U253/GND (-594 , 998)
*       104 = UAC36/U247/Gnd (-568.5 , 997)
*       104 = UAC36/U246/Gnd (-520.5 , 997)
*       104 = UAC37/U254/Gnd (-318 , 997)
*       104 = UAC37/U253/GND (-229.5 , 998)
*       104 = UAC37/U247/Gnd (-204 , 997)
*       104 = UAC37/U246/Gnd (-156 , 997)
*       104 = UAC38/U254/Gnd (45.5 , 997)
*       104 = UAC38/U253/GND (134 , 998)
*       104 = UAC38/U247/Gnd (159.5 , 997)
*       104 = UAC38/U246/Gnd (207.5 , 997)
*       104 = UAC112/U224/GND (-1921 , 1039.5)
*       104 = UAC112/U227/GND (-1799.5 , 1085)
*       104 = UAC112/U223/GND (-1866 , 1085)
*       104 = UAC112/U222/GND (-1883 , 1084.5)
*       104 = UAC112/U226/GND (-1837 , 1039.5)
*       104 = UAC112/U225/GND (-1854 , 1039)
*       104 = UAC112/U230/GND (-1753 , 1039.5)
*       104 = UAC112/U229/GND (-1770 , 1039)
*       104 = UAC112/U228/GND (-1774 , 1085)
*       104 = UAC78/U238/GND (-1497 , 1040.5)
*       104 = UAC78/U219/GND (-1496.5 , 1084.5)
*       104 = UAC78/U238/A (-1532 , 1053)
*       104 = UAC78/U219/A (-1531.5 , 1097)
*       104 = UAC78/U245/Gnd (-1474 , 1041)
*       104 = UAC78/U218/Gnd (-1447 , 1038)
*       104 = UAC78/U262/GND (-1475.5 , 1084.5)
*       104 = UAC78/U222/Gnd (-1453.5 , 1082)
*       104 = UAC78/U206/Gnd (-1323 , 1082)
*       104 = UAC78/U220/GND (-1325 , 1084.5)
*       104 = UAC78/U229/Gnd (-1340 , 1041)
*       104 = UAC78/U235/A (-1305.5 , 1053)
*       104 = UAC78/U236/GND (-1226 , 1040.5)
*       104 = UAC78/U235/GND (-1270.5 , 1040.5)
*       104 = UAC35/U262/GND (-1111.5 , 1084.5)
*       104 = UAC35/U245/Gnd (-1110 , 1041)
*       104 = UAC35/U238/GND (-1133 , 1040.5)
*       104 = UAC35/U219/GND (-1132.5 , 1084.5)
*       104 = UAC35/U218/Gnd (-1083 , 1038)
*       104 = UAC35/U222/Gnd (-1089.5 , 1082)
*       104 = UAC35/U206/Gnd (-959 , 1082)
*       104 = UAC35/U220/GND (-961 , 1084.5)
*       104 = UAC35/U235/GND (-906.5 , 1040.5)
*       104 = UAC35/U229/Gnd (-976 , 1041)
*       104 = UAC35/U236/GND (-862 , 1040.5)
*       104 = UAC36/U245/Gnd (-746.5 , 1041)
*       104 = UAC36/U238/GND (-769.5 , 1040.5)
*       104 = UAC36/U218/Gnd (-719.5 , 1038)
*       104 = UAC36/U262/GND (-748 , 1084.5)
*       104 = UAC36/U222/Gnd (-726 , 1082)
*       104 = UAC36/U219/GND (-769 , 1084.5)
*       104 = UAC36/U206/Gnd (-595.5 , 1082)
*       104 = UAC36/U220/GND (-597.5 , 1084.5)
*       104 = UAC36/U229/Gnd (-612.5 , 1041)
*       104 = UAC36/U236/GND (-498.5 , 1040.5)
*       104 = UAC36/U235/GND (-543 , 1040.5)
*       104 = UAC37/U238/GND (-405 , 1040.5)
*       104 = UAC37/U219/GND (-404.5 , 1084.5)
*       104 = UAC37/U245/Gnd (-382 , 1041)
*       104 = UAC37/U218/Gnd (-355 , 1038)
*       104 = UAC37/U262/GND (-383.5 , 1084.5)
*       104 = UAC37/U222/Gnd (-361.5 , 1082)
*       104 = UAC37/U206/Gnd (-231 , 1082)
*       104 = UAC37/U220/GND (-233 , 1084.5)
*       104 = UAC37/U229/Gnd (-248 , 1041)
*       104 = UAC37/U236/GND (-134 , 1040.5)
*       104 = UAC37/U235/GND (-178.5 , 1040.5)
*       104 = UAC38/U262/GND (-20 , 1084.5)
*       104 = UAC38/U222/Gnd (2 , 1082)
*       104 = UAC38/U219/GND (-41 , 1084.5)
*       104 = UAC38/U245/Gnd (-18.5 , 1041)
*       104 = UAC38/U238/GND (-41.5 , 1040.5)
*       104 = UAC38/U218/Gnd (8.5 , 1038)
*       104 = UAC38/U206/Gnd (132.5 , 1082)
*       104 = UAC38/U220/GND (130.5 , 1084.5)
*       104 = UAC38/U235/GND (185 , 1040.5)
*       104 = UAC38/U229/Gnd (115.5 , 1041)
*       104 = UAC38/U236/GND (229.5 , 1040.5)
*       104 = UAC38/U236/B (221 , 1053)
*       104 = UAC38/C (261.5 , 1080)
*       104 = UAC111/U224/GND (-1555.5 , 1202)
*       104 = UAC111/U232/GND (-1492.5 , 1157)
*       104 = UAC111/U231/GND (-1509.5 , 1156.5)
*       104 = UAC111/U229/GND (-1404.5 , 1201.5)
*       104 = UAC111/U226/GND (-1471.5 , 1202)
*       104 = UAC111/U225/GND (-1488.5 , 1201.5)
*       104 = UAC111/U220/Gnd (-1464 , 1154)
*       104 = UAC111/U230/GND (-1387.5 , 1202)
*       104 = UAC31/U245/Gnd (-1109.5 , 1203.5)
*       104 = UAC31/U238/GND (-1132.5 , 1203)
*       104 = UAC31/U254/Gnd (-1045.5 , 1159.5)
*       104 = UAC31/U218/Gnd (-1082.5 , 1200.5)
*       104 = UAC31/U235/GND (-906 , 1203)
*       104 = UAC31/U229/Gnd (-975.5 , 1203.5)
*       104 = UAC31/U253/GND (-957 , 1160.5)
*       104 = UAC31/U247/Gnd (-931.5 , 1159.5)
*       104 = UAC31/U236/GND (-861.5 , 1203)
*       104 = UAC31/U246/Gnd (-883.5 , 1159.5)
*       104 = UAC32/U245/Gnd (-746 , 1203.5)
*       104 = UAC32/U238/GND (-769 , 1203)
*       104 = UAC32/U218/Gnd (-719 , 1200.5)
*       104 = UAC32/U229/Gnd (-612 , 1203.5)
*       104 = UAC32/U254/Gnd (-682 , 1159.5)
*       104 = UAC32/U253/GND (-593.5 , 1160.5)
*       104 = UAC32/U236/GND (-498 , 1203)
*       104 = UAC32/U235/GND (-542.5 , 1203)
*       104 = UAC32/U247/Gnd (-568 , 1159.5)
*       104 = UAC32/U246/Gnd (-520 , 1159.5)
*       104 = UAC33/U238/GND (-404.5 , 1203)
*       104 = UAC33/U254/Gnd (-317.5 , 1159.5)
*       104 = UAC33/U245/Gnd (-381.5 , 1203.5)
*       104 = UAC33/U218/Gnd (-354.5 , 1200.5)
*       104 = UAC33/U229/Gnd (-247.5 , 1203.5)
*       104 = UAC33/U253/GND (-229 , 1160.5)
*       104 = UAC33/U247/Gnd (-203.5 , 1159.5)
*       104 = UAC33/U236/GND (-133.5 , 1203)
*       104 = UAC33/U235/GND (-178 , 1203)
*       104 = UAC33/U246/Gnd (-155.5 , 1159.5)
*       104 = UAC34/U245/Gnd (-18 , 1203.5)
*       104 = UAC34/U238/GND (-41 , 1203)
*       104 = UAC34/U218/Gnd (9 , 1200.5)
*       104 = UAC34/U254/Gnd (46 , 1159.5)
*       104 = UAC38/C6 (95.5 , 1129)
*       104 = UAC34/U235/GND (185.5 , 1203)
*       104 = UAC34/U229/Gnd (116 , 1203.5)
*       104 = UAC34/U253/GND (134.5 , 1160.5)
*       104 = UAC34/U247/Gnd (160 , 1159.5)
*       104 = UAC34/U246/Gnd (208 , 1159.5)
*       104 = UAC34/U236/GND (230 , 1203)
*       104 = UAC111/U223/GND (-1500.5 , 1247.5)
*       104 = UAC111/U222/GND (-1517.5 , 1247)
*       104 = UAC111/U228/GND (-1408.5 , 1247.5)
*       104 = UAC111/U227/GND (-1434 , 1247.5)
*       104 = UAC31/U262/GND (-1111 , 1247)
*       104 = UAC31/U219/GND (-1132 , 1247)
*       104 = UAC31/U222/Gnd (-1089 , 1244.5)
*       104 = UAC31/U206/Gnd (-958.5 , 1244.5)
*       104 = UAC31/U220/GND (-960.5 , 1247)
*       104 = UAC31/U206/A (-955 , 1264.5)
*       104 = UAC31/A6 (-953.5 , 1294)
*       104 = UAC32/U262/GND (-747.5 , 1247)
*       104 = UAC32/U222/Gnd (-725.5 , 1244.5)
*       104 = UAC32/U219/GND (-768.5 , 1247)
*       104 = UAC32/U206/Gnd (-595 , 1244.5)
*       104 = UAC32/U220/GND (-597 , 1247)
*       104 = UAC32/A6 (-590 , 1294)
*       104 = UAC33/U219/GND (-404 , 1247)
*       104 = UAC33/U262/GND (-383 , 1247)
*       104 = UAC33/U222/Gnd (-361 , 1244.5)
*       104 = UAC33/U206/Gnd (-230.5 , 1244.5)
*       104 = UAC33/U220/GND (-232.5 , 1247)
*       104 = UAC33/U206/A (-227 , 1264.5)
*       104 = UAC33/A6 (-225.5 , 1294)
*       104 = UAC33/U222/B (-284 , 1259.5)
*       104 = UAC34/U262/GND (-19.5 , 1247)
*       104 = UAC34/U222/Gnd (2.5 , 1244.5)
*       104 = UAC34/U219/GND (-40.5 , 1247)
*       104 = UAC34/U206/Gnd (133 , 1244.5)
*       104 = UAC34/U220/GND (131 , 1247)
*       104 = UAC34/U236/B (221.5 , 1215.5)
*       104 = UAC34/C (262 , 1242.5)
*       106 = UAC33/U246/Vin (-160.5 , 1173)
*       106 = UAC33/U236/OUT (-155 , 1204)
*       108 = UAC33/U253/B (-266 , 1162)
*       108 = UAC33/U246/Vout (-146.5 , 1173)
*       109 = UAC33/U253/C (-238.5 , 1161.5)
*       109 = UAC33/U247/Vout (-194.5 , 1173)
*       110 = UAC33/U247/Vin (-208.5 , 1173)
*       110 = UAC33/U235/OUT (-199.5 , 1204)
*       111 = UAC33/U229/Vin (-252.5 , 1217)
*       111 = UAC33/U220/OUT (-254 , 1248)
*       117 = UAC33/U245/Vout (-372.5 , 1217)
*       117 = UAC33/U253/A (-278.5 , 1161.5)
*       118 = UAC33/U254/Vin (-322.5 , 1173)
*       118 = UAC33/U253/OUT (-288 , 1161.5)
*       119 = UAC33/U218/A (-351 , 1220.5)
*       119 = UAC33/U222/Vout (-322 , 1271.5)
*       122 = UAC33/U238/OUT (-426 , 1204)
*       122 = UAC33/U245/Vin (-386.5 , 1217)
*       123 = UAC41/U219/A (-440 , 934.5)
*       123 = UAC37/B6 (-440 , 1024)
*       123 = UAC73/U238/A (-443.5 , -82.5)
*       123 = UAC73/B6 (-443.5 , -111.5)
*       123 = UAC73/U219/A (-443 , -38.5)
*       123 = UAC73/U235/A (-217 , -82.5)
*       123 = UAC69/U238/A (-443 , 80)
*       123 = UAC69/U219/A (-442.5 , 124)
*       123 = UAC69/B6 (-443 , 51)
*       123 = UAC69/U235/A (-216.5 , 80)
*       123 = UAC64/B6 (-442.5 , 212.5)
*       123 = UAC64/U238/A (-442.5 , 241.5)
*       123 = UAC64/U219/A (-442 , 285.5)
*       123 = UAC64/U235/A (-216 , 241.5)
*       123 = UAC60/U238/A (-442 , 404)
*       123 = UAC60/B6 (-442 , 375)
*       123 = UAC60/U235/A (-215.5 , 404)
*       123 = UAC60/U219/A (-441.5 , 448)
*       123 = UAC57/U238/A (-441.5 , 566.5)
*       123 = UAC57/U219/A (-441 , 610.5)
*       123 = UAC57/B6 (-441.5 , 537.5)
*       123 = UAC57/U235/A (-215 , 566.5)
*       123 = UAC53/B6 (-441 , 700)
*       123 = UAC53/U238/A (-441 , 729)
*       123 = UAC53/U219/A (-440.5 , 773)
*       123 = UAC53/U235/A (-214.5 , 729)
*       123 = UAC41/U238/A (-440.5 , 890.5)
*       123 = UAC41/B6 (-440.5 , 861.5)
*       123 = UAC41/U235/A (-214 , 890.5)
*       123 = UAC37/U238/A (-440 , 1053)
*       123 = UAC37/U219/A (-439.5 , 1097)
*       123 = UAC37/U235/A (-213.5 , 1053)
*       123 = UAC33/U238/A (-439.5 , 1215.5)
*       123 = UAC33/B6 (-439.5 , 1186.5)
*       123 = UAC33/U219/A (-439 , 1259.5)
*       123 = Bf1 (-439 , 1299)
*       123 = UAC33/U235/A (-213 , 1215.5)
*       124 = UAC33/U238/B (-413 , 1215.5)
*       124 = UAC33/U220/A (-267.5 , 1259.5)
*       124 = UAC33/C6 (-267.5 , 1291.5)
*       124 = UAC34/U254/Vout (55 , 1173)
*       124 = UAC34/P (56 , 1146)
*       124 = UAC33/U236/B (-142 , 1215.5)
*       124 = UAC33/C (-101.5 , 1242.5)
*       126 = UAC32/U247/Vin (-573 , 1173)
*       126 = UAC32/U235/OUT (-564 , 1204)
*       127 = UAC32/U246/Vin (-525 , 1173)
*       127 = UAC32/U236/OUT (-519.5 , 1204)
*       128 = UAC32/U236/A (-533 , 1215.5)
*       128 = UAC32/U235/B (-551 , 1215.5)
*       128 = UAC32/U206/Vout (-556 , 1271.5)
*       132 = UAC32/U218/B (-642 , 1215.5)
*       132 = UAC32/U229/Vout (-603 , 1217)
*       133 = UAC32/U254/Vin (-687 , 1173)
*       133 = UAC32/U253/OUT (-652.5 , 1161.5)
*       134 = UAC32/U253/B (-630.5 , 1162)
*       134 = UAC32/U246/Vout (-511 , 1173)
*       135 = UAC32/U253/C (-603 , 1161.5)
*       135 = UAC32/U247/Vout (-559 , 1173)
*       136 = UAC32/U229/Vin (-617 , 1217)
*       136 = UAC32/U220/OUT (-618.5 , 1248)
*       142 = UAC32/U245/Vout (-737 , 1217)
*       142 = UAC32/U253/A (-643 , 1161.5)
*       143 = UAC32/U218/A (-715.5 , 1220.5)
*       143 = UAC32/U222/Vout (-686.5 , 1271.5)
*       144 = UAC32/U245/Vin (-751 , 1217)
*       144 = UAC32/U238/OUT (-790.5 , 1204)
*       145 = UAC36/B6 (-804.5 , 1024)
*       145 = UAC40/U219/A (-804.5 , 934.5)
*       145 = UAC72/U238/A (-808 , -82.5)
*       145 = UAC72/B6 (-808 , -111.5)
*       145 = UAC72/U219/A (-807.5 , -38.5)
*       145 = UAC72/U235/A (-581.5 , -82.5)
*       145 = UAC68/U238/A (-807.5 , 80)
*       145 = UAC68/U219/A (-807 , 124)
*       145 = UAC68/B6 (-807.5 , 51)
*       145 = UAC68/U235/A (-581 , 80)
*       145 = UAC63/B6 (-807 , 212.5)
*       145 = UAC63/U238/A (-807 , 241.5)
*       145 = UAC63/U219/A (-806.5 , 285.5)
*       145 = UAC63/U235/A (-580.5 , 241.5)
*       145 = UAC66/U238/A (-806.5 , 404)
*       145 = UAC66/B6 (-806.5 , 375)
*       145 = UAC66/U235/A (-580 , 404)
*       145 = UAC66/U219/A (-806 , 448)
*       145 = UAC56/U238/A (-806 , 566.5)
*       145 = UAC56/U219/A (-805.5 , 610.5)
*       145 = UAC56/B6 (-806 , 537.5)
*       145 = UAC56/U235/A (-579.5 , 566.5)
*       145 = UAC52/B6 (-805.5 , 700)
*       145 = UAC52/U238/A (-805.5 , 729)
*       145 = UAC52/U219/A (-805 , 773)
*       145 = UAC52/U235/A (-579 , 729)
*       145 = UAC40/U238/A (-805 , 890.5)
*       145 = UAC40/B6 (-805 , 861.5)
*       145 = UAC40/U235/A (-578.5 , 890.5)
*       145 = UAC36/U238/A (-804.5 , 1053)
*       145 = UAC36/U219/A (-804 , 1097)
*       145 = UAC36/U235/A (-578 , 1053)
*       145 = UAC32/U238/A (-804 , 1215.5)
*       145 = UAC32/B6 (-804 , 1186.5)
*       145 = UAC32/U219/A (-803.5 , 1259.5)
*       145 = Bf2 (-803.5 , 1298)
*       145 = UAC32/U235/A (-577.5 , 1215.5)
*       146 = UAC31/U246/Vin (-888.5 , 1173)
*       146 = UAC31/U236/OUT (-883 , 1204)
*       148 = UAC32/U238/B (-777.5 , 1215.5)
*       148 = UAC32/U220/A (-632 , 1259.5)
*       148 = UAC32/C6 (-632 , 1291.5)
*       148 = UAC32/U236/B (-506.5 , 1215.5)
*       148 = UAC33/U254/Vout (-308.5 , 1173)
*       148 = UAC33/P (-307.5 , 1146)
*       148 = UAC32/C (-466 , 1242.5)
*       150 = UAC31/U253/C (-966.5 , 1161.5)
*       150 = UAC31/U247/Vout (-922.5 , 1173)
*       151 = UAC31/U247/Vin (-936.5 , 1173)
*       151 = UAC31/U235/OUT (-927.5 , 1204)
*       152 = UAC31/U236/A (-896.5 , 1215.5)
*       152 = UAC31/U235/B (-914.5 , 1215.5)
*       152 = UAC31/U206/Vout (-919.5 , 1271.5)
*       153 = UAC31/U229/Vin (-980.5 , 1217)
*       153 = UAC31/U220/OUT (-982 , 1248)
*       159 = UAC31/U218/B (-1005.5 , 1215.5)
*       159 = UAC31/U229/Vout (-966.5 , 1217)
*       160 = UAC31/U254/Vin (-1050.5 , 1173)
*       160 = UAC31/U253/OUT (-1016 , 1161.5)
*       161 = UAC31/U253/B (-994 , 1162)
*       161 = UAC31/U246/Vout (-874.5 , 1173)
*       162 = UAC31/U218/A (-1079 , 1220.5)
*       162 = UAC31/U222/Vout (-1050 , 1271.5)
*       165 = UAC31/U245/Vout (-1100.5 , 1217)
*       165 = UAC31/U253/A (-1006.5 , 1161.5)
*       166 = UAC31/U245/Vin (-1114.5 , 1217)
*       166 = UAC31/U238/OUT (-1154 , 1204)
*       167 = UAC39/U219/A (-1168 , 934.5)
*       167 = UAC35/B6 (-1168 , 1024)
*       167 = UAC71/U238/A (-1171.5 , -82.5)
*       167 = UAC71/B6 (-1171.5 , -111.5)
*       167 = UAC71/U219/A (-1171 , -38.5)
*       167 = UAC71/U235/A (-945 , -82.5)
*       167 = UAC67/U238/A (-1171 , 80)
*       167 = UAC67/U219/A (-1170.5 , 124)
*       167 = UAC67/B6 (-1171 , 51)
*       167 = UAC67/U235/A (-944.5 , 80)
*       167 = UAC62/B6 (-1170.5 , 212.5)
*       167 = UAC62/U238/A (-1170.5 , 241.5)
*       167 = UAC62/U219/A (-1170 , 285.5)
*       167 = UAC62/U235/A (-944 , 241.5)
*       167 = UAC59/U238/A (-1170 , 404)
*       167 = UAC59/B6 (-1170 , 375)
*       167 = UAC59/U235/A (-943.5 , 404)
*       167 = UAC59/U219/A (-1169.5 , 448)
*       167 = UAC55/U238/A (-1169.5 , 566.5)
*       167 = UAC55/U219/A (-1169 , 610.5)
*       167 = UAC55/B6 (-1169.5 , 537.5)
*       167 = UAC55/U235/A (-943 , 566.5)
*       167 = UAC51/B6 (-1169 , 700)
*       167 = UAC51/U238/A (-1169 , 729)
*       167 = UAC51/U219/A (-1168.5 , 773)
*       167 = UAC51/U235/A (-942.5 , 729)
*       167 = UAC39/U238/A (-1168.5 , 890.5)
*       167 = UAC39/B6 (-1168.5 , 861.5)
*       167 = UAC39/U235/A (-942 , 890.5)
*       167 = UAC35/U238/A (-1168 , 1053)
*       167 = UAC35/U219/A (-1167.5 , 1097)
*       167 = UAC35/U235/A (-941.5 , 1053)
*       167 = UAC31/U238/A (-1167.5 , 1215.5)
*       167 = UAC31/B6 (-1167.5 , 1186.5)
*       167 = UAC31/U219/A (-1167 , 1259.5)
*       167 = Bf3 (-1166.5 , 1298.5)
*       167 = UAC31/U235/A (-941 , 1215.5)
*       172 = UAC111/U230/vin (-1395.5 , 1214)
*       172 = UAC111/U229/OUT (-1426 , 1202.5)
*       173 = UAC111/U220/A (-1460.5 , 1174)
*       173 = UAC111/U232/vout (-1472 , 1168)
*       174 = UAC111/U226/vout (-1451 , 1213)
*       174 = UAC111/U227/B (-1445.5 , 1274)
*       179 = UAC111/U231/B (-1518 , 1169)
*       179 = UAC111/Pn (-1518.5 , 1142.5)
*       179 = UAC31/U254/Vout (-1036.5 , 1173)
*       179 = UAC31/P (-1035.5 , 1146)
*       180 = UAC111/U232/vin (-1500.5 , 1169)
*       180 = UAC111/U231/OUT (-1531 , 1157.5)
*       181 = UAC111/U225/OUT (-1510 , 1202.5)
*       181 = UAC111/U226/vin (-1479.5 , 1214)
*       182 = UAC111/U225/A (-1523.5 , 1214)
*       182 = UAC111/U224/vout (-1535 , 1213)
*       183 = UAC111/U225/B (-1497 , 1214)
*       183 = UAC111/U222/B (-1526 , 1259.5)
*       183 = UAC111/L (-1527 , 1297)
*       183 = Lf7 (-1526.5 , 1303.5)
*       186 = Q7 (-1803.5 , 1172)
*       186 = UAC112/Fn (-1956.5 , 1063)
*       186 = UAC112/U229/B (-1778.5 , 1051.5)
*       186 = UAC112/F (-1775 , 1137)
*       186 = UAC111/Qn (-1590.5 , 1172)
*       186 = UAC111/U220/Vout (-1425 , 1181)
*       190 = UAC38/U206/Vout (171.5 , 1109)
*       190 = UAC38/U236/A (194.5 , 1053)
*       190 = UAC38/U235/B (176.5 , 1053)
*       202 = UAC38/U218/B (85.5 , 1053)
*       202 = UAC38/U229/Vout (124.5 , 1054.5)
*       203 = UAC38/U222/Vout (41 , 1109)
*       203 = UAC38/U218/A (12 , 1058)
*       204 = UAC38/U229/Vin (110.5 , 1054.5)
*       204 = UAC38/U220/OUT (109 , 1085.5)
*       206 = UAC112/U228/vout (-1753.5 , 1096)
*       206 = UAC112/D (-1717 , 1091.5)
*       206 = UAC78/D (-1569.5 , 1093.5)
*       206 = UAC78/U219/B (-1505 , 1097)
*       206 = UAC78/D6 (-1505.5 , 1124)
*       206 = UAC78/U220/B (-1333.5 , 1097)
*       206 = UAC35/D (-1205.5 , 1093.5)
*       206 = UAC35/U219/B (-1141 , 1097)
*       206 = UAC35/D6 (-1141.5 , 1124)
*       206 = UAC35/U220/B (-969.5 , 1097)
*       206 = UAC36/D (-842 , 1093.5)
*       206 = UAC36/U219/B (-777.5 , 1097)
*       206 = UAC36/D6 (-778 , 1124)
*       206 = UAC36/U220/B (-606 , 1097)
*       206 = UAC37/D (-477.5 , 1093.5)
*       206 = UAC37/U219/B (-413 , 1097)
*       206 = UAC37/D6 (-413.5 , 1124)
*       206 = UAC37/U220/B (-241.5 , 1097)
*       206 = UAC38/D (-114 , 1093.5)
*       206 = UAC38/U219/B (-49.5 , 1097)
*       206 = UAC38/D6 (-50 , 1124)
*       206 = UAC38/U220/B (122 , 1097)
*       206 = UAC112/Dn (-1755 , 1138)
*       213 = UAC38/U219/OUT (-62.5 , 1085.5)
*       213 = UAC38/U262/vin (-12.5 , 1097.5)
*       214 = UAC38/U262/vout (-27 , 1099)
*       214 = UAC38/U222/A (5.5 , 1102)
*       215 = UAC38/U245/Vout (-9.5 , 1054.5)
*       215 = UAC38/U253/A (84.5 , 999)
*       216 = UAC38/U245/Vin (-23.5 , 1054.5)
*       216 = UAC38/U238/OUT (-63 , 1041.5)
*       223 = UAC37/U229/Vin (-253 , 1054.5)
*       223 = UAC37/U220/OUT (-254.5 , 1085.5)
*       227 = UAC37/U206/Vout (-192 , 1109)
*       227 = UAC37/U236/A (-169 , 1053)
*       227 = UAC37/U235/B (-187 , 1053)
*       235 = UAC37/U222/Vout (-322.5 , 1109)
*       235 = UAC37/U218/A (-351.5 , 1058)
*       238 = UAC37/U218/B (-278 , 1053)
*       238 = UAC37/U229/Vout (-239 , 1054.5)
*       244 = UAC37/U206/A (-227.5 , 1102)
*       244 = UAC37/U222/B (-284.5 , 1097)
*       244 = UAC37/A6 (-226 , 1131.5)
*       244 = UAC34/S (-117.5 , 1175.5)
*       244 = UAC34/U218/Vout (48 , 1227.5)
*       245 = UAC37/U219/OUT (-426 , 1085.5)
*       245 = UAC37/U262/vin (-376 , 1097.5)
*       246 = UAC37/U222/A (-358 , 1102)
*       246 = UAC37/U262/vout (-390.5 , 1099)
*       247 = UAC37/U238/B (-413.5 , 1053)
*       247 = UAC37/U220/A (-268 , 1097)
*       247 = UAC38/U254/Vout (54.5 , 1010.5)
*       247 = UAC38/P (55.5 , 983.5)
*       247 = UAC37/U236/B (-142.5 , 1053)
*       247 = UAC37/C (-102 , 1080)
*       247 = UAC37/C6 (-268 , 1129)
*       248 = UAC37/U238/OUT (-426.5 , 1041.5)
*       248 = UAC37/U245/Vin (-387 , 1054.5)
*       254 = UAC36/U206/Vout (-556.5 , 1109)
*       254 = UAC36/U236/A (-533.5 , 1053)
*       254 = UAC36/U235/B (-551.5 , 1053)
*       262 = UAC36/U206/A (-592 , 1102)
*       262 = UAC36/U222/B (-649 , 1097)
*       262 = UAC36/A6 (-590.5 , 1131.5)
*       262 = UAC33/S (-481 , 1175.5)
*       262 = UAC33/U218/Vout (-315.5 , 1227.5)
*       263 = UAC36/U218/B (-642.5 , 1053)
*       263 = UAC36/U229/Vout (-603.5 , 1054.5)
*       264 = UAC36/U229/Vin (-617.5 , 1054.5)
*       264 = UAC36/U220/OUT (-619 , 1085.5)
*       275 = UAC36/U262/vout (-755 , 1099)
*       275 = UAC36/U222/A (-722.5 , 1102)
*       276 = UAC36/U218/A (-716 , 1058)
*       276 = UAC36/U222/Vout (-687 , 1109)
*       278 = UAC36/U219/OUT (-790.5 , 1085.5)
*       278 = UAC36/U262/vin (-740.5 , 1097.5)
*       279 = UAC36/U245/Vin (-751.5 , 1054.5)
*       279 = UAC36/U238/OUT (-791 , 1041.5)
*       282 = UAC36/U238/B (-778 , 1053)
*       282 = UAC36/U220/A (-632.5 , 1097)
*       282 = UAC36/U236/B (-507 , 1053)
*       282 = UAC37/U254/Vout (-309 , 1010.5)
*       282 = UAC37/P (-308 , 983.5)
*       282 = UAC36/C (-466.5 , 1080)
*       282 = UAC36/C6 (-632.5 , 1129)
*       287 = UAC35/U206/Vout (-920 , 1109)
*       287 = UAC35/U236/A (-897 , 1053)
*       287 = UAC35/U235/B (-915 , 1053)
*       288 = UAC35/U229/Vin (-981 , 1054.5)
*       288 = UAC35/U220/OUT (-982.5 , 1085.5)
*       300 = UAC35/U238/B (-1141.5 , 1053)
*       300 = UAC35/U220/A (-996 , 1097)
*       300 = UAC36/U254/Vout (-673.5 , 1010.5)
*       300 = UAC36/P (-672.5 , 983.5)
*       300 = UAC35/U236/B (-870.5 , 1053)
*       300 = UAC35/C (-830 , 1080)
*       300 = UAC35/C6 (-996 , 1129)
*       301 = UAC35/U222/B (-1012.5 , 1097)
*       301 = UAC35/U206/A (-955.5 , 1102)
*       301 = UAC35/A6 (-954 , 1131.5)
*       301 = UAC32/S (-845.5 , 1175.5)
*       301 = UAC32/U218/Vout (-680 , 1227.5)
*       302 = UAC35/U218/B (-1006 , 1053)
*       302 = UAC35/U229/Vout (-967 , 1054.5)
*       303 = UAC35/U222/Vout (-1050.5 , 1109)
*       303 = UAC35/U218/A (-1079.5 , 1058)
*       310 = UAC35/U219/OUT (-1154 , 1085.5)
*       310 = UAC35/U262/vin (-1104 , 1097.5)
*       311 = UAC35/U262/vout (-1118.5 , 1099)
*       311 = UAC35/U222/A (-1086 , 1102)
*       312 = UAC35/U245/Vout (-1101 , 1054.5)
*       312 = UAC35/U253/A (-1007 , 999)
*       313 = UAC35/U245/Vin (-1115 , 1054.5)
*       313 = UAC35/U238/OUT (-1154.5 , 1041.5)
*       323 = UAC78/U229/Vin (-1345 , 1054.5)
*       323 = UAC78/U220/OUT (-1346.5 , 1085.5)
*       325 = UAC78/U206/Vout (-1284 , 1109)
*       325 = UAC78/U236/A (-1261 , 1053)
*       325 = UAC78/U235/B (-1279 , 1053)
*       331 = UAC78/U262/vout (-1482.5 , 1099)
*       331 = UAC78/U222/A (-1450 , 1102)
*       332 = UAC78/U222/Vout (-1414.5 , 1109)
*       332 = UAC78/U218/A (-1443.5 , 1058)
*       333 = UAC78/U218/Vout (-1408 , 1065)
*       333 = UAC80/U222/B (-1740.5 , 934.5)
*       333 = UAC80/U206/A (-1683.5 , 939.5)
*       333 = UAC80/A6 (-1682 , 969)
*       333 = UAC78/S (-1573.5 , 1013)
*       335 = UAC78/U218/B (-1370 , 1053)
*       335 = UAC78/U229/Vout (-1331 , 1054.5)
*       337 = UAC78/U206/A (-1319.5 , 1102)
*       337 = UAC78/U222/B (-1376.5 , 1097)
*       337 = UAC78/A6 (-1318 , 1131.5)
*       337 = UAC31/S (-1209 , 1175.5)
*       337 = UAC31/U218/Vout (-1043.5 , 1227.5)
*       344 = UAC78/U219/OUT (-1518 , 1085.5)
*       344 = UAC78/U262/vin (-1468 , 1097.5)
*       345 = UAC78/U238/B (-1505.5 , 1053)
*       345 = UAC78/U220/A (-1360 , 1097)
*       345 = UAC35/U254/Vout (-1037 , 1010.5)
*       345 = UAC35/P (-1036 , 983.5)
*       345 = UAC78/U236/B (-1234.5 , 1053)
*       345 = UAC78/C (-1194 , 1080)
*       345 = UAC78/C6 (-1360 , 1129)
*       346 = UAC78/U238/OUT (-1518.5 , 1041.5)
*       346 = UAC78/U245/Vin (-1479 , 1054.5)
*       349 = UAC112/U229/OUT (-1791.5 , 1040)
*       349 = UAC112/U230/vin (-1761 , 1051.5)
*       350 = UAC112/U226/vin (-1845 , 1051.5)
*       350 = UAC112/U225/OUT (-1875.5 , 1040)
*       351 = UAC112/U227/B (-1811 , 1111.5)
*       351 = UAC112/U226/vout (-1816.5 , 1050.5)
*       352 = UAC112/U227/O/P (-1797.5 , 1105)
*       352 = UAC112/U228/vin (-1782 , 1097)
*       353 = UAC112/U223/vout (-1845.5 , 1096)
*       353 = UAC112/An (-1846.5 , 1140)
*       353 = UAC38/U222/B (79 , 1097)
*       353 = UAC38/U206/A (136 , 1102)
*       353 = UAC38/A6 (137.5 , 1131.5)
*       357 = UAC112/U222/B (-1891.5 , 1097)
*       357 = UAC112/U225/B (-1862.5 , 1051.5)
*       357 = UAC112/L (-1892.5 , 1134.5)
*       357 = Lf6 (-1892 , 1139)
*       358 = UAC112/U222/OUT (-1904.5 , 1085.5)
*       358 = UAC112/U223/vin (-1874 , 1097)
*       359 = UAC112/U224/vout (-1900.5 , 1050.5)
*       359 = UAC112/U225/A (-1889 , 1051.5)
*       363 = UAC38/U246/Vin (202.5 , 1010.5)
*       363 = UAC38/U236/OUT (208 , 1041.5)
*       364 = UAC38/U253/C (124.5 , 999)
*       364 = UAC38/U247/Vout (168.5 , 1010.5)
*       365 = UAC38/U247/Vin (154.5 , 1010.5)
*       365 = UAC38/U235/OUT (163.5 , 1041.5)
*       371 = UAC38/U253/B (97 , 999.5)
*       371 = UAC38/U246/Vout (216.5 , 1010.5)
*       372 = UAC38/U254/Vin (40.5 , 1010.5)
*       372 = UAC38/U253/OUT (75 , 999)
*       380 = UAC37/U246/Vin (-161 , 1010.5)
*       380 = UAC37/U236/OUT (-155.5 , 1041.5)
*       384 = UAC37/U253/B (-266.5 , 999.5)
*       384 = UAC37/U246/Vout (-147 , 1010.5)
*       385 = UAC37/U253/C (-239 , 999)
*       385 = UAC37/U247/Vout (-195 , 1010.5)
*       386 = UAC37/U247/Vin (-209 , 1010.5)
*       386 = UAC37/U235/OUT (-200 , 1041.5)
*       391 = UAC41/U206/Vout (-192.5 , 946.5)
*       391 = UAC41/U236/A (-169.5 , 890.5)
*       391 = UAC41/U235/B (-187.5 , 890.5)
*       395 = UAC37/U245/Vout (-373 , 1054.5)
*       395 = UAC37/U253/A (-279 , 999)
*       396 = UAC37/U254/Vin (-323 , 1010.5)
*       396 = UAC37/U253/OUT (-288.5 , 999)
*       400 = UAC41/U206/A (-228 , 939.5)
*       400 = UAC41/A6 (-226.5 , 969)
*       400 = UAC41/U222/B (-285 , 934.5)
*       400 = UAC38/S (-118 , 1013)
*       400 = UAC38/U218/Vout (47.5 , 1065)
*       404 = UAC36/U247/Vin (-573.5 , 1010.5)
*       404 = UAC36/U235/OUT (-564.5 , 1041.5)
*       405 = UAC36/U246/Vin (-525.5 , 1010.5)
*       405 = UAC36/U236/OUT (-520 , 1041.5)
*       409 = UAC36/U254/Vin (-687.5 , 1010.5)
*       409 = UAC36/U253/OUT (-653 , 999)
*       410 = UAC36/U253/B (-631 , 999.5)
*       410 = UAC36/U246/Vout (-511.5 , 1010.5)
*       411 = UAC36/U253/C (-603.5 , 999)
*       411 = UAC36/U247/Vout (-559.5 , 1010.5)
*       419 = UAC36/U245/Vout (-737.5 , 1054.5)
*       419 = UAC36/U253/A (-643.5 , 999)
*       422 = UAC35/U246/Vin (-889 , 1010.5)
*       422 = UAC35/U236/OUT (-883.5 , 1041.5)
*       426 = UAC35/U253/C (-967 , 999)
*       426 = UAC35/U247/Vout (-923 , 1010.5)
*       427 = UAC35/U247/Vin (-937 , 1010.5)
*       427 = UAC35/U235/OUT (-928 , 1041.5)
*       430 = UAC114/U220/B (-2129.5 , 844)
*       430 = UAC114/U230/vout (-2109.5 , 888)
*       430 = UAC114/Fn (-2093.5 , 912)
*       430 = UAC80/F (-1933.5 , 943)
*       430 = UAC80/U206/B (-1610 , 934.5)
*       430 = UAC80/F6 (-1606 , 963)
*       430 = UAC79/F (-1570 , 943)
*       430 = UAC79/U206/B (-1246.5 , 934.5)
*       430 = UAC79/F6 (-1242.5 , 963)
*       430 = UAC39/F (-1206 , 943)
*       430 = UAC40/F (-842.5 , 943)
*       430 = UAC39/U206/B (-882.5 , 934.5)
*       430 = UAC39/F6 (-878.5 , 963)
*       430 = UAC40/U206/B (-519 , 934.5)
*       430 = UAC40/F6 (-515 , 963)
*       430 = UAC41/F (-478 , 943)
*       430 = UAC42/F (-114.5 , 943)
*       430 = UAC41/U206/B (-154.5 , 934.5)
*       430 = UAC41/F6 (-150.5 , 963)
*       430 = UAC42/U206/B (209 , 934.5)
*       430 = UAC42/F6 (213 , 963)
*       436 = UAC35/U254/Vin (-1051 , 1010.5)
*       436 = UAC35/U253/OUT (-1016.5 , 999)
*       437 = UAC35/U253/B (-994.5 , 999.5)
*       437 = UAC35/U246/Vout (-875 , 1010.5)
*       443 = UAC78/U246/Vin (-1253 , 1010.5)
*       443 = UAC78/U236/OUT (-1247.5 , 1041.5)
*       449 = UAC78/U253/B (-1358.5 , 999.5)
*       449 = UAC78/U246/Vout (-1239 , 1010.5)
*       450 = UAC78/U253/C (-1331 , 999)
*       450 = UAC78/U247/Vout (-1287 , 1010.5)
*       451 = UAC78/U247/Vin (-1301 , 1010.5)
*       451 = UAC78/U235/OUT (-1292 , 1041.5)
*       457 = UAC78/U245/Vout (-1465 , 1054.5)
*       457 = UAC78/U253/A (-1371 , 999)
*       458 = UAC78/U254/Vin (-1415 , 1010.5)
*       458 = UAC78/U253/OUT (-1380.5 , 999)
*       460 = UAC79/U206/A (-1320 , 939.5)
*       460 = UAC79/A6 (-1318.5 , 969)
*       460 = UAC79/U222/B (-1377 , 934.5)
*       460 = UAC35/S (-1209.5 , 1013)
*       460 = UAC35/U218/Vout (-1044 , 1065)
*       469 = UAC112/U220/B (-1752.5 , 1006.5)
*       469 = UAC112/U230/vout (-1732.5 , 1050.5)
*       469 = UAC112/Fn (-1716.5 , 1074.5)
*       469 = UAC78/F (-1569.5 , 1105.5)
*       469 = UAC78/U206/B (-1246 , 1097)
*       469 = UAC35/F (-1205.5 , 1105.5)
*       469 = UAC78/F6 (-1242 , 1125.5)
*       469 = UAC36/F (-842 , 1105.5)
*       469 = UAC35/U206/B (-882 , 1097)
*       469 = UAC35/F6 (-878 , 1125.5)
*       469 = UAC36/U206/B (-518.5 , 1097)
*       469 = UAC37/F (-477.5 , 1105.5)
*       469 = UAC36/F6 (-514.5 , 1125.5)
*       469 = UAC38/F (-114 , 1105.5)
*       469 = UAC37/U206/B (-154 , 1097)
*       469 = UAC37/F6 (-150 , 1125.5)
*       469 = UAC38/U206/B (209.5 , 1097)
*       469 = UAC38/F6 (213.5 , 1125.5)
*       480 = UAC112/U220/A (-1826 , 1011.5)
*       480 = UAC112/U232/vout (-1837.5 , 1005.5)
*       482 = UAC114/Fn (-2333.5 , 900.5)
*       482 = UAC114/U229/B (-2155.5 , 889)
*       482 = UAC114/F (-2152 , 974.5)
*       482 = Q6 (-2179 , 1009.5)
*       482 = UAC112/Qn (-1956 , 1009.5)
*       482 = UAC112/U220/Vout (-1790.5 , 1018.5)
*       485 = UAC112/U231/OUT (-1896.5 , 995)
*       485 = UAC112/U232/vin (-1866 , 1006.5)
*       487 = UAC112/U231/B (-1883.5 , 1006.5)
*       487 = UAC112/Pn (-1884 , 980)
*       487 = UAC78/U254/Vout (-1401 , 1010.5)
*       487 = UAC78/P (-1400 , 983.5)
*       489 = UAC114/U228/vin (-2159 , 934.5)
*       489 = UAC114/U227/O/P (-2174.5 , 942.5)
*       491 = UAC125/B (-1280.5 , -38.5)
*       491 = UAC121/U224/vin (-4093.5 , 78.5)
*       491 = UAC121/Z (-4119 , 112)
*       491 = UAC121/U231/A (-4074.5 , 33.5)
*       491 = UAC121/U222/A (-4082.5 , 124)
*       491 = UAC121/U229/A (-3969.5 , 78.5)
*       491 = UAC121/U227/A (-3991 , 140)
*       491 = UAC120/Z (-3808 , 273.5)
*       491 = UAC120/U231/A (-3763.5 , 195)
*       491 = UAC120/U224/vin (-3782.5 , 240)
*       491 = UAC120/U222/A (-3771.5 , 285.5)
*       491 = UAC120/U229/A (-3658.5 , 240)
*       491 = UAC120/U227/A (-3680 , 301.5)
*       491 = UAC119/U231/A (-3398.5 , 357.5)
*       491 = UAC119/U224/vin (-3417.5 , 402.5)
*       491 = UAC119/U222/A (-3406.5 , 448)
*       491 = UAC119/Z (-3443 , 436)
*       491 = UAC119/U229/A (-3293.5 , 402.5)
*       491 = UAC119/U227/A (-3315 , 464)
*       491 = UAC118/U231/A (-3024 , 520)
*       491 = UAC118/U224/vin (-3043 , 565)
*       491 = UAC118/U222/A (-3032 , 610.5)
*       491 = UAC118/Z (-3068.5 , 598.5)
*       491 = UAC118/U229/A (-2919 , 565)
*       491 = UAC118/U227/A (-2940.5 , 626.5)
*       491 = UAC116/Z (-2702.5 , 761)
*       491 = UAC116/U231/A (-2658 , 682.5)
*       491 = UAC116/U224/vin (-2677 , 727.5)
*       491 = UAC116/U222/A (-2666 , 773)
*       491 = UAC116/U229/A (-2553 , 727.5)
*       491 = UAC116/U227/A (-2574.5 , 789)
*       491 = UAC114/U224/vin (-2306 , 889)
*       491 = UAC114/Z (-2331.5 , 922.5)
*       491 = UAC114/U231/A (-2287 , 844)
*       491 = UAC114/U222/A (-2295 , 934.5)
*       491 = UAC114/U227/A (-2203.5 , 950.5)
*       491 = UAC114/U229/A (-2182 , 889)
*       491 = UAC112/U231/A (-1910 , 1006.5)
*       491 = UAC112/U224/vin (-1929 , 1051.5)
*       491 = UAC112/U222/A (-1918 , 1097)
*       491 = UAC112/Z (-1954.5 , 1085)
*       491 = UAC112/U229/A (-1805 , 1051.5)
*       491 = UAC112/U227/A (-1826.5 , 1113)
*       491 = UAC111/U231/A (-1544.5 , 1169)
*       491 = UAC111/U224/vin (-1563.5 , 1214)
*       491 = UAC111/U222/A (-1552.5 , 1259.5)
*       491 = UAC111/Z (-1589 , 1247.5)
*       491 = UAC111/U229/A (-1439.5 , 1214)
*       491 = UAC111/U227/A (-1461 , 1275.5)
*       493 = UAC42/U253/C (124 , 836.5)
*       493 = UAC42/U247/Vout (168 , 848)
*       494 = UAC42/U236/A (194 , 890.5)
*       494 = UAC42/U235/B (176 , 890.5)
*       494 = UAC42/U206/Vout (171 , 946.5)
*       495 = UAC42/U247/Vin (154 , 848)
*       495 = UAC42/U235/OUT (163 , 879)
*       498 = UAC42/U246/Vin (202 , 848)
*       498 = UAC42/U236/OUT (207.5 , 879)
*       503 = UAC42/U220/B (121.5 , 934.5)
*       503 = UAC42/U219/B (-50 , 934.5)
*       503 = UAC42/D6 (-50.5 , 961.5)
*       503 = UAC41/U220/B (-242 , 934.5)
*       503 = UAC40/U220/B (-606.5 , 934.5)
*       503 = UAC40/U219/B (-778 , 934.5)
*       503 = UAC40/D6 (-778.5 , 961.5)
*       503 = UAC39/U220/B (-970 , 934.5)
*       503 = UAC79/U220/B (-1334 , 934.5)
*       503 = UAC80/U220/B (-1697.5 , 934.5)
*       503 = UAC80/U219/B (-1869 , 934.5)
*       503 = UAC80/D6 (-1869.5 , 961.5)
*       503 = UAC114/U228/vout (-2130.5 , 933.5)
*       503 = UAC114/D (-2094 , 929)
*       503 = UAC114/Dn (-2132 , 975.5)
*       503 = UAC80/D (-1933.5 , 931)
*       503 = UAC79/D (-1570 , 931)
*       503 = UAC79/U219/B (-1505.5 , 934.5)
*       503 = UAC79/D6 (-1506 , 961.5)
*       503 = UAC39/D (-1206 , 931)
*       503 = UAC39/U219/B (-1141.5 , 934.5)
*       503 = UAC39/D6 (-1142 , 961.5)
*       503 = UAC40/D (-842.5 , 931)
*       503 = UAC41/D (-478 , 931)
*       503 = UAC41/U219/B (-413.5 , 934.5)
*       503 = UAC41/D6 (-414 , 961.5)
*       503 = UAC42/D (-114.5 , 931)
*       504 = UAC42/U218/B (85 , 890.5)
*       504 = UAC42/U229/Vout (124 , 892)
*       505 = UAC42/U253/B (96.5 , 837)
*       505 = UAC42/U246/Vout (216 , 848)
*       506 = UAC42/U222/B (78.5 , 934.5)
*       506 = UAC114/U223/vout (-2222.5 , 933.5)
*       506 = UAC114/An (-2223.5 , 977.5)
*       506 = UAC42/U206/A (135.5 , 939.5)
*       506 = UAC42/A6 (137 , 969)
*       507 = UAC42/U218/A (11.5 , 895.5)
*       507 = UAC42/U222/Vout (40.5 , 946.5)
*       508 = UAC42/U220/OUT (108.5 , 923)
*       508 = UAC42/U229/Vin (110 , 892)
*       510 = UAC42/U254/Vin (40 , 848)
*       510 = UAC42/U253/OUT (74.5 , 836.5)
*       515 = UAC42/U262/vin (-13 , 935)
*       515 = UAC42/U219/OUT (-63 , 923)
*       516 = UAC42/U245/Vout (-10 , 892)
*       516 = UAC42/U253/A (84 , 836.5)
*       517 = UAC42/U245/Vin (-24 , 892)
*       517 = UAC42/U238/OUT (-63.5 , 879)
*       518 = UAC42/U262/vout (-27.5 , 936.5)
*       518 = UAC42/U222/A (5 , 939.5)
*       520 = UAC41/U246/Vin (-161.5 , 848)
*       520 = UAC41/U236/OUT (-156 , 879)
*       523 = UAC41/U253/B (-267 , 837)
*       523 = UAC41/U246/Vout (-147.5 , 848)
*       524 = UAC41/U253/C (-239.5 , 836.5)
*       524 = UAC41/U247/Vout (-195.5 , 848)
*       525 = UAC41/U247/Vin (-209.5 , 848)
*       525 = UAC41/U235/OUT (-200.5 , 879)
*       526 = UAC41/U229/Vin (-253.5 , 892)
*       526 = UAC41/U220/OUT (-255 , 923)
*       533 = UAC41/U245/Vout (-373.5 , 892)
*       533 = UAC41/U253/A (-279.5 , 836.5)
*       534 = UAC41/U254/Vin (-323.5 , 848)
*       534 = UAC41/U253/OUT (-289 , 836.5)
*       535 = UAC41/U218/A (-352 , 895.5)
*       535 = UAC41/U222/Vout (-323 , 946.5)
*       538 = UAC41/U218/B (-278.5 , 890.5)
*       538 = UAC41/U229/Vout (-239.5 , 892)
*       541 = UAC41/U238/OUT (-427 , 879)
*       541 = UAC41/U245/Vin (-387.5 , 892)
*       542 = UAC41/U222/A (-358.5 , 939.5)
*       542 = UAC41/U262/vout (-391 , 936.5)
*       543 = UAC41/U238/B (-414 , 890.5)
*       543 = UAC41/U220/A (-268.5 , 934.5)
*       543 = UAC41/C6 (-268.5 , 966.5)
*       543 = UAC42/P (55 , 821)
*       543 = UAC41/U236/B (-143 , 890.5)
*       543 = UAC41/C (-102.5 , 917.5)
*       543 = UAC42/U254/Vout (54 , 848)
*       544 = UAC41/U219/OUT (-426.5 , 923)
*       544 = UAC41/U262/vin (-376.5 , 935)
*       547 = UAC40/U236/A (-534 , 890.5)
*       547 = UAC40/U235/B (-552 , 890.5)
*       547 = UAC40/U206/Vout (-557 , 946.5)
*       548 = UAC40/U247/Vin (-574 , 848)
*       548 = UAC40/U235/OUT (-565 , 879)
*       549 = UAC40/U246/Vin (-526 , 848)
*       549 = UAC40/U236/OUT (-520.5 , 879)
*       553 = UAC40/U218/B (-643 , 890.5)
*       553 = UAC40/U229/Vout (-604 , 892)
*       554 = UAC40/U254/Vin (-688 , 848)
*       554 = UAC40/U253/OUT (-653.5 , 836.5)
*       555 = UAC40/U253/B (-631.5 , 837)
*       555 = UAC40/U246/Vout (-512 , 848)
*       556 = UAC40/U253/C (-604 , 836.5)
*       556 = UAC40/U247/Vout (-560 , 848)
*       557 = UAC40/U229/Vin (-618 , 892)
*       557 = UAC40/U220/OUT (-619.5 , 923)
*       558 = UAC40/U206/A (-592.5 , 939.5)
*       558 = UAC40/U222/B (-649.5 , 934.5)
*       558 = UAC40/A6 (-591 , 969)
*       558 = UAC37/S (-481.5 , 1013)
*       558 = UAC37/U218/Vout (-316 , 1065)
*       566 = UAC40/U262/vin (-741 , 935)
*       566 = UAC40/U219/OUT (-791 , 923)
*       567 = UAC40/U245/Vout (-738 , 892)
*       567 = UAC40/U253/A (-644 , 836.5)
*       568 = UAC40/U262/vout (-755.5 , 936.5)
*       568 = UAC40/U222/A (-723 , 939.5)
*       569 = UAC40/U218/A (-716.5 , 895.5)
*       569 = UAC40/U222/Vout (-687.5 , 946.5)
*       570 = UAC40/U238/OUT (-791.5 , 879)
*       570 = UAC40/U245/Vin (-752 , 892)
*       571 = UAC39/U246/Vin (-889.5 , 848)
*       571 = UAC39/U236/OUT (-884 , 879)
*       573 = UAC40/U238/B (-778.5 , 890.5)
*       573 = UAC40/U220/A (-633 , 934.5)
*       573 = UAC40/C6 (-633 , 966.5)
*       573 = UAC40/U236/B (-507.5 , 890.5)
*       573 = UAC41/P (-308.5 , 821)
*       573 = UAC40/C (-467 , 917.5)
*       573 = UAC41/U254/Vout (-309.5 , 848)
*       576 = UAC39/U253/C (-967.5 , 836.5)
*       576 = UAC39/U247/Vout (-923.5 , 848)
*       577 = UAC39/U236/A (-897.5 , 890.5)
*       577 = UAC39/U235/B (-915.5 , 890.5)
*       577 = UAC39/U206/Vout (-920.5 , 946.5)
*       578 = UAC39/U247/Vin (-937.5 , 848)
*       578 = UAC39/U235/OUT (-928.5 , 879)
*       579 = UAC39/U229/Vin (-981.5 , 892)
*       579 = UAC39/U220/OUT (-983 , 923)
*       586 = UAC39/U218/B (-1006.5 , 890.5)
*       586 = UAC39/U229/Vout (-967.5 , 892)
*       587 = UAC39/U254/Vin (-1051.5 , 848)
*       587 = UAC39/U253/OUT (-1017 , 836.5)
*       588 = UAC39/U253/B (-995 , 837)
*       588 = UAC39/U246/Vout (-875.5 , 848)
*       589 = UAC39/U222/B (-1013 , 934.5)
*       589 = UAC39/U206/A (-956 , 939.5)
*       589 = UAC39/A6 (-954.5 , 969)
*       589 = UAC36/S (-846 , 1013)
*       589 = UAC36/U218/Vout (-680.5 , 1065)
*       590 = UAC39/U218/A (-1080 , 895.5)
*       590 = UAC39/U222/Vout (-1051 , 946.5)
*       595 = UAC39/U262/vin (-1104.5 , 935)
*       595 = UAC39/U219/OUT (-1154.5 , 923)
*       596 = UAC39/U245/Vout (-1101.5 , 892)
*       596 = UAC39/U253/A (-1007.5 , 836.5)
*       597 = UAC39/U245/Vin (-1115.5 , 892)
*       597 = UAC39/U238/OUT (-1155 , 879)
*       598 = UAC39/U262/vout (-1119 , 936.5)
*       598 = UAC39/U222/A (-1086.5 , 939.5)
*       599 = UAC39/U238/B (-1142 , 890.5)
*       599 = UAC39/U220/A (-996.5 , 934.5)
*       599 = UAC39/C6 (-996.5 , 966.5)
*       599 = UAC40/P (-673 , 821)
*       599 = UAC39/U236/B (-871 , 890.5)
*       599 = UAC39/C (-830.5 , 917.5)
*       599 = UAC40/U254/Vout (-674 , 848)
*       602 = UAC79/U246/Vin (-1253.5 , 848)
*       602 = UAC79/U236/OUT (-1248 , 879)
*       604 = UAC79/U253/B (-1359 , 837)
*       604 = UAC79/U246/Vout (-1239.5 , 848)
*       605 = UAC79/U253/C (-1331.5 , 836.5)
*       605 = UAC79/U247/Vout (-1287.5 , 848)
*       606 = UAC79/U247/Vin (-1301.5 , 848)
*       606 = UAC79/U235/OUT (-1292.5 , 879)
*       607 = UAC79/U229/Vin (-1345.5 , 892)
*       607 = UAC79/U220/OUT (-1347 , 923)
*       608 = UAC79/U236/A (-1261.5 , 890.5)
*       608 = UAC79/U235/B (-1279.5 , 890.5)
*       608 = UAC79/U206/Vout (-1284.5 , 946.5)
*       615 = UAC79/U245/Vout (-1465.5 , 892)
*       615 = UAC79/U253/A (-1371.5 , 836.5)
*       616 = UAC79/U254/Vin (-1415.5 , 848)
*       616 = UAC79/U253/OUT (-1381 , 836.5)
*       617 = UAC79/U262/vout (-1483 , 936.5)
*       617 = UAC79/U222/A (-1450.5 , 939.5)
*       618 = UAC79/U218/A (-1444 , 895.5)
*       618 = UAC79/U222/Vout (-1415 , 946.5)
*       620 = UAC79/U218/B (-1370.5 , 890.5)
*       620 = UAC79/U229/Vout (-1331.5 , 892)
*       624 = UAC79/U238/OUT (-1519 , 879)
*       624 = UAC79/U245/Vin (-1479.5 , 892)
*       625 = UAC79/U238/B (-1506 , 890.5)
*       625 = UAC79/U220/A (-1360.5 , 934.5)
*       625 = UAC79/C6 (-1360.5 , 966.5)
*       625 = UAC39/P (-1036.5 , 821)
*       625 = UAC79/U236/B (-1235 , 890.5)
*       625 = UAC79/C (-1194.5 , 917.5)
*       625 = UAC39/U254/Vout (-1037.5 , 848)
*       626 = UAC79/U219/OUT (-1518.5 , 923)
*       626 = UAC79/U262/vin (-1468.5 , 935)
*       629 = UAC80/U236/A (-1625 , 890.5)
*       629 = UAC80/U235/B (-1643 , 890.5)
*       629 = UAC80/U206/Vout (-1648 , 946.5)
*       630 = UAC80/U247/Vin (-1665 , 848)
*       630 = UAC80/U235/OUT (-1656 , 879)
*       631 = UAC80/U246/Vin (-1617 , 848)
*       631 = UAC80/U236/OUT (-1611.5 , 879)
*       637 = UAC80/U218/B (-1734 , 890.5)
*       637 = UAC80/U229/Vout (-1695 , 892)
*       638 = UAC80/U254/Vin (-1779 , 848)
*       638 = UAC80/U253/OUT (-1744.5 , 836.5)
*       639 = UAC80/U253/B (-1722.5 , 837)
*       639 = UAC80/U246/Vout (-1603 , 848)
*       640 = UAC80/U253/C (-1695 , 836.5)
*       640 = UAC80/U247/Vout (-1651 , 848)
*       641 = UAC80/U229/Vin (-1709 , 892)
*       641 = UAC80/U220/OUT (-1710.5 , 923)
*       648 = UAC80/U262/vin (-1832 , 935)
*       648 = UAC80/U219/OUT (-1882 , 923)
*       649 = UAC80/U245/Vout (-1829 , 892)
*       649 = UAC80/U253/A (-1735 , 836.5)
*       650 = UAC80/U245/Vin (-1843 , 892)
*       650 = UAC80/U238/OUT (-1882.5 , 879)
*       651 = UAC80/U238/B (-1869.5 , 890.5)
*       651 = UAC80/U220/A (-1724 , 934.5)
*       651 = UAC80/C6 (-1724 , 966.5)
*       651 = UAC80/U236/B (-1598.5 , 890.5)
*       651 = UAC79/P (-1400.5 , 821)
*       651 = UAC80/C (-1558 , 917.5)
*       651 = UAC79/U254/Vout (-1401.5 , 848)
*       652 = UAC80/U262/vout (-1846.5 , 936.5)
*       652 = UAC80/U222/A (-1814 , 939.5)
*       653 = UAC80/U218/A (-1807.5 , 895.5)
*       653 = UAC80/U222/Vout (-1778.5 , 946.5)
*       657 = UAC114/U227/B (-2188 , 949)
*       657 = UAC114/U226/vout (-2193.5 , 888)
*       658 = UAC114/U230/vin (-2138 , 889)
*       658 = UAC114/U229/OUT (-2168.5 , 877.5)
*       664 = UAC114/U222/B (-2268.5 , 934.5)
*       664 = UAC114/L (-2269.5 , 972)
*       664 = Lf5 (-2269.5 , 977)
*       664 = UAC114/U225/B (-2239.5 , 889)
*       665 = UAC114/U232/vin (-2243 , 844)
*       665 = UAC114/U231/OUT (-2273.5 , 832.5)
*       666 = UAC114/U226/vin (-2222 , 889)
*       666 = UAC114/U225/OUT (-2252.5 , 877.5)
*       667 = UAC114/U222/OUT (-2281.5 , 923)
*       667 = UAC114/U223/vin (-2251 , 934.5)
*       668 = UAC114/U220/A (-2203 , 849)
*       668 = UAC114/U232/vout (-2214.5 , 843)
*       671 = UAC114/U225/A (-2266 , 889)
*       671 = UAC114/U224/vout (-2277.5 , 888)
*       681 = UAC54/U222/B (78 , 773)
*       681 = UAC116/U223/vout (-2593.5 , 772)
*       681 = UAC116/An (-2594.5 , 816)
*       681 = UAC54/U206/A (135 , 778)
*       681 = UAC54/A6 (136.5 , 807.5)
*       682 = UAC54/U220/OUT (108 , 761.5)
*       682 = UAC54/U229/Vin (109.5 , 730.5)
*       683 = UAC116/U228/vout (-2501.5 , 772)
*       683 = UAC116/Dn (-2503 , 814)
*       683 = UAC116/D (-2465 , 767.5)
*       683 = UAC84/D (-2310 , 769.5)
*       683 = UAC84/U219/B (-2245.5 , 773)
*       683 = UAC84/D6 (-2246 , 800)
*       683 = UAC84/U220/B (-2074 , 773)
*       683 = UAC82/D (-1946.5 , 769.5)
*       683 = UAC82/U219/B (-1882 , 773)
*       683 = UAC82/D6 (-1882.5 , 800)
*       683 = UAC82/U220/B (-1710.5 , 773)
*       683 = UAC81/D (-1578 , 769.5)
*       683 = UAC81/U219/B (-1513.5 , 773)
*       683 = UAC81/D6 (-1514 , 800)
*       683 = UAC81/U220/B (-1342 , 773)
*       683 = UAC51/D (-1206.5 , 769.5)
*       683 = UAC51/U219/B (-1142 , 773)
*       683 = UAC51/D6 (-1142.5 , 800)
*       683 = UAC51/U220/B (-970.5 , 773)
*       683 = UAC52/D (-843 , 769.5)
*       683 = UAC52/U219/B (-778.5 , 773)
*       683 = UAC52/D6 (-779 , 800)
*       683 = UAC52/U220/B (-607 , 773)
*       683 = UAC53/D (-478.5 , 769.5)
*       683 = UAC53/U219/B (-414 , 773)
*       683 = UAC53/D6 (-414.5 , 800)
*       683 = UAC53/U220/B (-242.5 , 773)
*       683 = UAC54/D (-115 , 769.5)
*       683 = UAC54/U219/B (-50.5 , 773)
*       683 = UAC54/D6 (-51 , 800)
*       683 = UAC54/U220/B (121 , 773)
*       690 = UAC54/U219/OUT (-63.5 , 761.5)
*       690 = UAC54/U262/vin (-13.5 , 773.5)
*       691 = UAC54/U262/vout (-28 , 775)
*       691 = UAC54/U222/A (4.5 , 778)
*       698 = UAC53/U206/Vout (-193 , 785)
*       698 = UAC53/U236/A (-170 , 729)
*       698 = UAC53/U235/B (-188 , 729)
*       710 = UAC53/U206/A (-228.5 , 778)
*       710 = UAC53/A6 (-227 , 807.5)
*       710 = UAC53/U222/B (-285.5 , 773)
*       710 = UAC42/S (-118.5 , 850.5)
*       710 = UAC42/U218/Vout (47 , 902.5)
*       711 = UAC53/U219/OUT (-427 , 761.5)
*       711 = UAC53/U262/vin (-377 , 773.5)
*       712 = UAC53/U262/vout (-391.5 , 775)
*       712 = UAC53/U222/A (-359 , 778)
*       720 = UAC52/U206/A (-593 , 778)
*       720 = UAC52/A6 (-591.5 , 807.5)
*       720 = UAC52/U222/B (-650 , 773)
*       720 = UAC41/S (-482 , 850.5)
*       720 = UAC41/U218/Vout (-316.5 , 902.5)
*       728 = UAC52/U262/vout (-756 , 775)
*       728 = UAC52/U222/A (-723.5 , 778)
*       731 = UAC52/U219/OUT (-791.5 , 761.5)
*       731 = UAC52/U262/vin (-741.5 , 773.5)
*       738 = UAC116/U220/B (-2500.5 , 682.5)
*       738 = UAC116/U230/vout (-2480.5 , 726.5)
*       738 = UAC116/Fn (-2464.5 , 750.5)
*       738 = UAC84/F (-2310 , 781.5)
*       738 = UAC84/U206/B (-1986.5 , 773)
*       738 = UAC84/F6 (-1982.5 , 801.5)
*       738 = UAC82/F (-1946.5 , 781.5)
*       738 = UAC82/U206/B (-1623 , 773)
*       738 = UAC82/F6 (-1619 , 801.5)
*       738 = UAC81/F (-1578 , 781.5)
*       738 = UAC81/U206/B (-1254.5 , 773)
*       738 = UAC81/F6 (-1250.5 , 801.5)
*       738 = UAC51/F (-1206.5 , 781.5)
*       738 = UAC52/F (-843 , 781.5)
*       738 = UAC51/U206/B (-883 , 773)
*       738 = UAC51/F6 (-879 , 801.5)
*       738 = UAC52/U206/B (-519.5 , 773)
*       738 = UAC52/F6 (-515.5 , 801.5)
*       738 = UAC53/F (-478.5 , 781.5)
*       738 = UAC54/F (-115 , 781.5)
*       738 = UAC53/U206/B (-155 , 773)
*       738 = UAC53/F6 (-151 , 801.5)
*       738 = UAC54/U206/B (208.5 , 773)
*       738 = UAC54/F6 (212.5 , 801.5)
*       744 = UAC51/U222/B (-1013.5 , 773)
*       744 = UAC51/U206/A (-956.5 , 778)
*       744 = UAC51/A6 (-955 , 807.5)
*       744 = UAC40/S (-846.5 , 850.5)
*       744 = UAC40/U218/Vout (-681 , 902.5)
*       750 = UAC51/U219/OUT (-1155 , 761.5)
*       750 = UAC51/U262/vin (-1105 , 773.5)
*       751 = UAC51/U262/vout (-1119.5 , 775)
*       751 = UAC51/U222/A (-1087 , 778)
*       758 = UAC81/U206/Vout (-1292.5 , 785)
*       758 = UAC81/U236/A (-1269.5 , 729)
*       758 = UAC81/U235/B (-1287.5 , 729)
*       770 = UAC81/U206/A (-1328 , 778)
*       770 = UAC81/A6 (-1326.5 , 807.5)
*       770 = UAC81/U222/B (-1385 , 773)
*       770 = UAC39/S (-1210 , 850.5)
*       770 = UAC39/U218/Vout (-1044.5 , 902.5)
*       771 = UAC81/U219/OUT (-1526.5 , 761.5)
*       771 = UAC81/U262/vin (-1476.5 , 773.5)
*       772 = UAC81/U222/A (-1458.5 , 778)
*       772 = UAC81/U262/vout (-1491 , 775)
*       780 = UAC82/U206/A (-1696.5 , 778)
*       780 = UAC82/A6 (-1695 , 807.5)
*       780 = UAC82/U222/B (-1753.5 , 773)
*       780 = UAC79/S (-1574 , 850.5)
*       780 = UAC79/U218/Vout (-1408.5 , 902.5)
*       787 = UAC82/U262/vout (-1859.5 , 775)
*       787 = UAC82/U222/A (-1827 , 778)
*       789 = UAC82/U218/A (-1820.5 , 734)
*       789 = UAC82/U222/Vout (-1791.5 , 785)
*       792 = UAC82/U219/OUT (-1895 , 761.5)
*       792 = UAC82/U262/vin (-1845 , 773.5)
*       799 = UAC84/U246/Vin (-1993.5 , 686.5)
*       799 = UAC84/U236/OUT (-1988 , 717.5)
*       805 = UAC84/U222/B (-2117 , 773)
*       805 = UAC84/U206/A (-2060 , 778)
*       805 = UAC84/A6 (-2058.5 , 807.5)
*       805 = UAC80/S (-1937.5 , 850.5)
*       805 = UAC80/U218/Vout (-1772 , 902.5)
*       811 = UAC114/Pn (-2261 , 817.5)
*       811 = UAC114/U231/B (-2260.5 , 844)
*       811 = UAC80/P (-1764 , 821)
*       811 = UAC80/U254/Vout (-1765 , 848)
*       812 = UAC84/U219/OUT (-2258.5 , 761.5)
*       812 = UAC84/U262/vin (-2208.5 , 773.5)
*       813 = UAC84/U262/vout (-2223 , 775)
*       813 = UAC84/U222/A (-2190.5 , 778)
*       815 = UAC116/U228/vin (-2530 , 773)
*       815 = UAC116/U227/O/P (-2545.5 , 781)
*       817 = UAC116/U223/vin (-2622 , 773)
*       817 = UAC116/U222/OUT (-2652.5 , 761.5)
*       819 = UAC116/Fn (-2704.5 , 739)
*       819 = UAC116/U229/B (-2526.5 , 727.5)
*       819 = UAC116/F (-2523 , 813)
*       819 = Q5 (-2549 , 846.5)
*       819 = UAC114/Qn (-2333 , 847)
*       819 = UAC114/U220/Vout (-2167.5 , 856)
*       820 = UAC54/U253/C (123.5 , 675)
*       820 = UAC54/U247/Vout (167.5 , 686.5)
*       821 = UAC54/U247/Vin (153.5 , 686.5)
*       821 = UAC54/U235/OUT (162.5 , 717.5)
*       822 = UAC54/U246/Vin (201.5 , 686.5)
*       822 = UAC54/U236/OUT (207 , 717.5)
*       824 = UAC54/U206/Vout (170.5 , 785)
*       824 = UAC54/U236/A (193.5 , 729)
*       824 = UAC54/U235/B (175.5 , 729)
*       828 = UAC54/U253/B (96 , 675.5)
*       828 = UAC54/U246/Vout (215.5 , 686.5)
*       829 = UAC54/U218/B (84.5 , 729)
*       829 = UAC54/U229/Vout (123.5 , 730.5)
*       830 = UAC54/U222/Vout (40 , 785)
*       830 = UAC54/U218/A (11 , 734)
*       833 = UAC54/U254/Vin (39.5 , 686.5)
*       833 = UAC54/U253/OUT (74 , 675)
*       836 = UAC54/U253/A (83.5 , 675)
*       836 = UAC54/U245/Vout (-10.5 , 730.5)
*       838 = UAC54/U238/OUT (-64 , 717.5)
*       838 = UAC54/U245/Vin (-24.5 , 730.5)
*       839 = UAC53/U246/Vin (-162 , 686.5)
*       839 = UAC53/U236/OUT (-156.5 , 717.5)
*       841 = UAC53/U253/B (-267.5 , 675.5)
*       841 = UAC53/U246/Vout (-148 , 686.5)
*       842 = UAC53/U253/C (-240 , 675)
*       842 = UAC53/U247/Vout (-196 , 686.5)
*       843 = UAC53/U247/Vin (-210 , 686.5)
*       843 = UAC53/U235/OUT (-201 , 717.5)
*       844 = UAC53/U229/Vin (-254 , 730.5)
*       844 = UAC53/U220/OUT (-255.5 , 761.5)
*       849 = UAC53/U253/A (-280 , 675)
*       849 = UAC53/U245/Vout (-374 , 730.5)
*       850 = UAC53/U254/Vin (-324 , 686.5)
*       850 = UAC53/U253/OUT (-289.5 , 675)
*       851 = UAC53/U229/Vout (-240 , 730.5)
*       851 = UAC53/U218/B (-279 , 729)
*       852 = UAC53/U222/Vout (-323.5 , 785)
*       852 = UAC53/U218/A (-352.5 , 734)
*       855 = UAC53/U238/OUT (-427.5 , 717.5)
*       855 = UAC53/U245/Vin (-388 , 730.5)
*       856 = UAC53/U238/B (-414.5 , 729)
*       856 = UAC53/U220/A (-269 , 773)
*       856 = UAC53/C6 (-269 , 805)
*       856 = UAC54/U254/Vout (53.5 , 686.5)
*       856 = UAC54/P (54.5 , 659.5)
*       856 = UAC53/U236/B (-143.5 , 729)
*       856 = UAC53/C (-103 , 756)
*       858 = UAC52/U247/Vin (-574.5 , 686.5)
*       858 = UAC52/U235/OUT (-565.5 , 717.5)
*       859 = UAC52/U246/Vin (-526.5 , 686.5)
*       859 = UAC52/U236/OUT (-521 , 717.5)
*       861 = UAC52/U206/Vout (-557.5 , 785)
*       861 = UAC52/U236/A (-534.5 , 729)
*       861 = UAC52/U235/B (-552.5 , 729)
*       864 = UAC52/U254/Vin (-688.5 , 686.5)
*       864 = UAC52/U253/OUT (-654 , 675)
*       865 = UAC52/U253/B (-632 , 675.5)
*       865 = UAC52/U246/Vout (-512.5 , 686.5)
*       866 = UAC52/U253/C (-604.5 , 675)
*       866 = UAC52/U247/Vout (-560.5 , 686.5)
*       867 = UAC52/U229/Vout (-604.5 , 730.5)
*       867 = UAC52/U218/B (-643.5 , 729)
*       869 = UAC52/U229/Vin (-618.5 , 730.5)
*       869 = UAC52/U220/OUT (-620 , 761.5)
*       874 = UAC52/U253/A (-644.5 , 675)
*       874 = UAC52/U245/Vout (-738.5 , 730.5)
*       875 = UAC52/U218/A (-717 , 734)
*       875 = UAC52/U222/Vout (-688 , 785)
*       876 = UAC52/U238/OUT (-792 , 717.5)
*       876 = UAC52/U245/Vin (-752.5 , 730.5)
*       877 = UAC51/U246/Vin (-890 , 686.5)
*       877 = UAC51/U236/OUT (-884.5 , 717.5)
*       879 = UAC52/U238/B (-779 , 729)
*       879 = UAC52/U220/A (-633.5 , 773)
*       879 = UAC52/C6 (-633.5 , 805)
*       879 = UAC52/U236/B (-508 , 729)
*       879 = UAC53/U254/Vout (-310 , 686.5)
*       879 = UAC53/P (-309 , 659.5)
*       879 = UAC52/C (-467.5 , 756)
*       881 = UAC51/U253/C (-968 , 675)
*       881 = UAC51/U247/Vout (-924 , 686.5)
*       882 = UAC51/U247/Vin (-938 , 686.5)
*       882 = UAC51/U235/OUT (-929 , 717.5)
*       883 = UAC51/U229/Vin (-982 , 730.5)
*       883 = UAC51/U220/OUT (-983.5 , 761.5)
*       885 = UAC51/U206/Vout (-921 , 785)
*       885 = UAC51/U236/A (-898 , 729)
*       885 = UAC51/U235/B (-916 , 729)
*       889 = UAC51/U254/Vin (-1052 , 686.5)
*       889 = UAC51/U253/OUT (-1017.5 , 675)
*       890 = UAC51/U218/B (-1007 , 729)
*       890 = UAC51/U229/Vout (-968 , 730.5)
*       891 = UAC51/U222/Vout (-1051.5 , 785)
*       891 = UAC51/U218/A (-1080.5 , 734)
*       894 = UAC51/U253/B (-995.5 , 675.5)
*       894 = UAC51/U246/Vout (-876 , 686.5)
*       896 = UAC51/U253/A (-1008 , 675)
*       896 = UAC51/U245/Vout (-1102 , 730.5)
*       897 = UAC51/U238/B (-1142.5 , 729)
*       897 = UAC51/U220/A (-997 , 773)
*       897 = UAC51/C6 (-997 , 805)
*       897 = UAC52/U254/Vout (-674.5 , 686.5)
*       897 = UAC52/P (-673.5 , 659.5)
*       897 = UAC51/U236/B (-871.5 , 729)
*       897 = UAC51/C (-831 , 756)
*       899 = UAC51/U238/OUT (-1155.5 , 717.5)
*       899 = UAC51/U245/Vin (-1116 , 730.5)
*       900 = UAC81/U246/Vin (-1261.5 , 686.5)
*       900 = UAC81/U236/OUT (-1256 , 717.5)
*       902 = UAC81/U253/B (-1367 , 675.5)
*       902 = UAC81/U246/Vout (-1247.5 , 686.5)
*       903 = UAC81/U253/C (-1339.5 , 675)
*       903 = UAC81/U247/Vout (-1295.5 , 686.5)
*       904 = UAC81/U247/Vin (-1309.5 , 686.5)
*       904 = UAC81/U235/OUT (-1300.5 , 717.5)
*       905 = UAC81/U229/Vin (-1353.5 , 730.5)
*       905 = UAC81/U220/OUT (-1355 , 761.5)
*       910 = UAC81/U253/A (-1379.5 , 675)
*       910 = UAC81/U245/Vout (-1473.5 , 730.5)
*       911 = UAC81/U254/Vin (-1423.5 , 686.5)
*       911 = UAC81/U253/OUT (-1389 , 675)
*       912 = UAC81/U229/Vout (-1339.5 , 730.5)
*       912 = UAC81/U218/B (-1378.5 , 729)
*       913 = UAC81/U222/Vout (-1423 , 785)
*       913 = UAC81/U218/A (-1452 , 734)
*       916 = UAC81/U238/OUT (-1527 , 717.5)
*       916 = UAC81/U245/Vin (-1487.5 , 730.5)
*       917 = UAC81/U238/B (-1514 , 729)
*       917 = UAC81/U220/A (-1368.5 , 773)
*       917 = UAC81/C6 (-1368.5 , 805)
*       917 = UAC51/U254/Vout (-1038 , 686.5)
*       917 = UAC51/P (-1037 , 659.5)
*       917 = UAC81/U236/B (-1243 , 729)
*       917 = UAC81/C (-1202.5 , 756)
*       919 = UAC82/U247/Vin (-1678 , 686.5)
*       919 = UAC82/U235/OUT (-1669 , 717.5)
*       920 = UAC82/U246/Vin (-1630 , 686.5)
*       920 = UAC82/U236/OUT (-1624.5 , 717.5)
*       922 = UAC82/U206/Vout (-1661 , 785)
*       922 = UAC82/U236/A (-1638 , 729)
*       922 = UAC82/U235/B (-1656 , 729)
*       925 = UAC82/U253/B (-1735.5 , 675.5)
*       925 = UAC82/U246/Vout (-1616 , 686.5)
*       926 = UAC82/U253/C (-1708 , 675)
*       926 = UAC82/U247/Vout (-1664 , 686.5)
*       927 = UAC82/U229/Vout (-1708 , 730.5)
*       927 = UAC82/U218/B (-1747 , 729)
*       929 = UAC82/U229/Vin (-1722 , 730.5)
*       929 = UAC82/U220/OUT (-1723.5 , 761.5)
*       934 = UAC82/U253/A (-1748 , 675)
*       934 = UAC82/U245/Vout (-1842 , 730.5)
*       935 = UAC82/U254/Vin (-1792 , 686.5)
*       935 = UAC82/U253/OUT (-1757.5 , 675)
*       936 = UAC82/U238/OUT (-1895.5 , 717.5)
*       936 = UAC82/U245/Vin (-1856 , 730.5)
*       937 = UAC82/U238/B (-1882.5 , 729)
*       937 = UAC82/U220/A (-1737 , 773)
*       937 = UAC82/C6 (-1737 , 805)
*       937 = UAC82/U236/B (-1611.5 , 729)
*       937 = UAC81/U254/Vout (-1409.5 , 686.5)
*       937 = UAC81/P (-1408.5 , 659.5)
*       937 = UAC82/C (-1571 , 756)
*       939 = UAC84/U253/C (-2071.5 , 675)
*       939 = UAC84/U247/Vout (-2027.5 , 686.5)
*       940 = UAC84/U247/Vin (-2041.5 , 686.5)
*       940 = UAC84/U235/OUT (-2032.5 , 717.5)
*       941 = UAC84/U229/Vin (-2085.5 , 730.5)
*       941 = UAC84/U220/OUT (-2087 , 761.5)
*       944 = UAC84/U206/Vout (-2024.5 , 785)
*       944 = UAC84/U236/A (-2001.5 , 729)
*       944 = UAC84/U235/B (-2019.5 , 729)
*       948 = UAC84/U254/Vin (-2155.5 , 686.5)
*       948 = UAC84/U253/OUT (-2121 , 675)
*       949 = UAC84/U253/B (-2099 , 675.5)
*       949 = UAC84/U246/Vout (-1979.5 , 686.5)
*       950 = UAC84/U218/B (-2110.5 , 729)
*       950 = UAC84/U229/Vout (-2071.5 , 730.5)
*       951 = UAC84/U222/Vout (-2155 , 785)
*       951 = UAC84/U218/A (-2184 , 734)
*       955 = UAC84/U253/A (-2111.5 , 675)
*       955 = UAC84/U245/Vout (-2205.5 , 730.5)
*       956 = UAC84/U238/B (-2246 , 729)
*       956 = UAC84/U220/A (-2100.5 , 773)
*       956 = UAC84/C6 (-2100.5 , 805)
*       956 = UAC82/U254/Vout (-1778 , 686.5)
*       956 = UAC82/P (-1777 , 659.5)
*       956 = UAC84/U236/B (-1975 , 729)
*       956 = UAC84/C (-1934.5 , 756)
*       958 = UAC84/U238/OUT (-2259 , 717.5)
*       958 = UAC84/U245/Vin (-2219.5 , 730.5)
*       962 = UAC116/U227/B (-2559 , 787.5)
*       962 = UAC116/U226/vout (-2564.5 , 726.5)
*       964 = UAC116/U229/OUT (-2539.5 , 716)
*       964 = UAC116/U230/vin (-2509 , 727.5)
*       968 = UAC116/U220/A (-2574 , 687.5)
*       968 = UAC116/U232/vout (-2585.5 , 681.5)
*       969 = UAC116/U231/B (-2631.5 , 682.5)
*       969 = UAC116/Pn (-2632 , 656)
*       969 = UAC84/U254/Vout (-2141.5 , 686.5)
*       969 = UAC84/P (-2140.5 , 659.5)
*       970 = UAC116/U232/vin (-2614 , 682.5)
*       970 = UAC116/U231/OUT (-2644.5 , 671)
*       971 = UAC116/U225/OUT (-2623.5 , 716)
*       971 = UAC116/U226/vin (-2593 , 727.5)
*       972 = UAC116/U225/A (-2637 , 727.5)
*       972 = UAC116/U224/vout (-2648.5 , 726.5)
*       973 = UAC116/U225/B (-2610.5 , 727.5)
*       973 = UAC116/U222/B (-2639.5 , 773)
*       973 = UAC116/L (-2640.5 , 810.5)
*       973 = Lf4 (-2640 , 815.5)
*       976 = Q4 (-2935.5 , 686)
*       976 = UAC118/Fn (-3070.5 , 576.5)
*       976 = UAC118/U229/B (-2892.5 , 565)
*       976 = UAC118/F (-2889 , 650.5)
*       976 = UAC116/Qn (-2704 , 685.5)
*       976 = UAC116/U220/Vout (-2538.5 , 694.5)
*       980 = UAC58/U206/Vout (170 , 622.5)
*       980 = UAC58/U236/A (193 , 566.5)
*       980 = UAC58/U235/B (175 , 566.5)
*       992 = UAC58/U218/B (84 , 566.5)
*       992 = UAC58/U229/Vout (123 , 568)
*       993 = UAC58/U220/OUT (107.5 , 599)
*       993 = UAC58/U229/Vin (109 , 568)
*       994 = UAC58/U222/B (77.5 , 610.5)
*       994 = UAC118/U223/vout (-2959.5 , 609.5)
*       994 = UAC118/An (-2960.5 , 653.5)
*       994 = UAC58/U206/A (134.5 , 615.5)
*       994 = UAC58/A6 (136 , 645)
*       995 = UAC58/U222/Vout (39.5 , 622.5)
*       995 = UAC58/U218/A (10.5 , 571.5)
*       997 = UAC118/U228/vout (-2867.5 , 609.5)
*       997 = UAC118/D (-2831 , 605)
*       997 = UAC90/D (-2681 , 607)
*       997 = UAC90/U219/B (-2616.5 , 610.5)
*       997 = UAC90/U220/B (-2445 , 610.5)
*       997 = UAC88/D (-2310.5 , 607)
*       997 = UAC88/U219/B (-2246 , 610.5)
*       997 = UAC88/U220/B (-2074.5 , 610.5)
*       997 = UAC87/D (-1946.5 , 607)
*       997 = UAC87/U219/B (-1882 , 610.5)
*       997 = UAC87/U220/B (-1710.5 , 610.5)
*       997 = UAC85/D (-1578.5 , 607)
*       997 = UAC85/U219/B (-1514 , 610.5)
*       997 = UAC85/U220/B (-1342.5 , 610.5)
*       997 = UAC55/D (-1207 , 607)
*       997 = UAC55/U219/B (-1142.5 , 610.5)
*       997 = UAC55/U220/B (-971 , 610.5)
*       997 = UAC56/D (-843.5 , 607)
*       997 = UAC56/U219/B (-779 , 610.5)
*       997 = UAC56/U220/B (-607.5 , 610.5)
*       997 = UAC57/D (-479 , 607)
*       997 = UAC57/U219/B (-414.5 , 610.5)
*       997 = UAC57/U220/B (-243 , 610.5)
*       997 = UAC58/D (-115.5 , 607)
*       997 = UAC58/U219/B (-51 , 610.5)
*       997 = UAC58/U220/B (120.5 , 610.5)
*       997 = UAC118/Dn (-2869 , 651.5)
*       997 = UAC90/D6 (-2617 , 637.5)
*       997 = UAC88/D6 (-2246.5 , 637.5)
*       997 = UAC87/D6 (-1882.5 , 637.5)
*       997 = UAC85/D6 (-1514.5 , 637.5)
*       997 = UAC55/D6 (-1143 , 637.5)
*       997 = UAC56/D6 (-779.5 , 637.5)
*       997 = UAC57/D6 (-415 , 637.5)
*       997 = UAC58/D6 (-51.5 , 637.5)
*       1006 = UAC58/U262/vout (-28.5 , 612.5)
*       1006 = UAC58/U222/A (4 , 615.5)
*       1007 = UAC58/U245/Vout (-11 , 568)
*       1007 = UAC58/U253/A (83 , 512.5)
*       1008 = UAC58/U245/Vin (-25 , 568)
*       1008 = UAC58/U238/OUT (-64.5 , 555)
*       1009 = UAC58/U262/vin (-14 , 611)
*       1009 = UAC58/U219/OUT (-64 , 599)
*       1015 = UAC57/U229/Vin (-254.5 , 568)
*       1015 = UAC57/U220/OUT (-256 , 599)
*       1022 = UAC57/U206/Vout (-193.5 , 622.5)
*       1022 = UAC57/U236/A (-170.5 , 566.5)
*       1022 = UAC57/U235/B (-188.5 , 566.5)
*       1031 = UAC57/U245/Vout (-374.5 , 568)
*       1031 = UAC57/U253/A (-280.5 , 512.5)
*       1032 = UAC57/U222/Vout (-324 , 622.5)
*       1032 = UAC57/U218/A (-353 , 571.5)
*       1034 = UAC57/U218/B (-279.5 , 566.5)
*       1034 = UAC57/U229/Vout (-240.5 , 568)
*       1040 = UAC57/U222/B (-286 , 610.5)
*       1040 = UAC57/U206/A (-229 , 615.5)
*       1040 = UAC57/A6 (-227.5 , 645)
*       1040 = UAC54/S (-119 , 689)
*       1040 = UAC54/U218/Vout (46.5 , 741)
*       1041 = UAC57/U262/vout (-392 , 612.5)
*       1041 = UAC57/U222/A (-359.5 , 615.5)
*       1042 = UAC57/U238/B (-415 , 566.5)
*       1042 = UAC57/U220/A (-269.5 , 610.5)
*       1042 = UAC58/U254/Vout (53 , 524)
*       1042 = UAC58/P (54 , 497)
*       1042 = UAC57/U236/B (-144 , 566.5)
*       1042 = UAC57/C (-103.5 , 593.5)
*       1042 = UAC57/C6 (-269.5 , 642.5)
*       1043 = UAC57/U238/OUT (-428 , 555)
*       1043 = UAC57/U245/Vin (-388.5 , 568)
*       1044 = UAC57/U219/OUT (-427.5 , 599)
*       1044 = UAC57/U262/vin (-377.5 , 611)
*       1050 = UAC56/U206/Vout (-558 , 622.5)
*       1050 = UAC56/U236/A (-535 , 566.5)
*       1050 = UAC56/U235/B (-553 , 566.5)
*       1057 = UAC56/U218/B (-644 , 566.5)
*       1057 = UAC56/U229/Vout (-605 , 568)
*       1058 = UAC56/U229/Vin (-619 , 568)
*       1058 = UAC56/U220/OUT (-620.5 , 599)
*       1059 = UAC56/U222/B (-650.5 , 610.5)
*       1059 = UAC56/U206/A (-593.5 , 615.5)
*       1059 = UAC56/A6 (-592 , 645)
*       1059 = UAC53/S (-482.5 , 689)
*       1059 = UAC53/U218/Vout (-317 , 741)
*       1072 = UAC56/U262/vout (-756.5 , 612.5)
*       1072 = UAC56/U222/A (-724 , 615.5)
*       1073 = UAC56/U245/Vout (-739 , 568)
*       1073 = UAC56/U253/A (-645 , 512.5)
*       1074 = UAC56/U218/A (-717.5 , 571.5)
*       1074 = UAC56/U222/Vout (-688.5 , 622.5)
*       1077 = UAC56/U238/OUT (-792.5 , 555)
*       1077 = UAC56/U245/Vin (-753 , 568)
*       1078 = UAC56/U219/OUT (-792 , 599)
*       1078 = UAC56/U262/vin (-742 , 611)
*       1081 = UAC56/U238/B (-779.5 , 566.5)
*       1081 = UAC56/U220/A (-634 , 610.5)
*       1081 = UAC56/U236/B (-508.5 , 566.5)
*       1081 = UAC57/U254/Vout (-310.5 , 524)
*       1081 = UAC57/P (-309.5 , 497)
*       1081 = UAC56/C (-468 , 593.5)
*       1081 = UAC56/C6 (-634 , 642.5)
*       1086 = UAC55/U206/Vout (-921.5 , 622.5)
*       1086 = UAC55/U236/A (-898.5 , 566.5)
*       1086 = UAC55/U235/B (-916.5 , 566.5)
*       1087 = UAC55/U229/Vin (-982.5 , 568)
*       1087 = UAC55/U220/OUT (-984 , 599)
*       1093 = UAC118/U220/B (-2866.5 , 520)
*       1093 = UAC118/U230/vout (-2846.5 , 564)
*       1093 = UAC118/Fn (-2830.5 , 588)
*       1093 = UAC90/F (-2681 , 619)
*       1093 = UAC90/U206/B (-2357.5 , 610.5)
*       1093 = UAC88/F (-2310.5 , 619)
*       1093 = UAC90/F6 (-2353.5 , 639)
*       1093 = UAC88/U206/B (-1987 , 610.5)
*       1093 = UAC87/F (-1946.5 , 619)
*       1093 = UAC88/F6 (-1983 , 639)
*       1093 = UAC87/U206/B (-1623 , 610.5)
*       1093 = UAC85/F (-1578.5 , 619)
*       1093 = UAC87/F6 (-1619 , 639)
*       1093 = UAC85/U206/B (-1255 , 610.5)
*       1093 = UAC55/F (-1207 , 619)
*       1093 = UAC85/F6 (-1251 , 639)
*       1093 = UAC56/F (-843.5 , 619)
*       1093 = UAC55/U206/B (-883.5 , 610.5)
*       1093 = UAC55/F6 (-879.5 , 639)
*       1093 = UAC56/U206/B (-520 , 610.5)
*       1093 = UAC57/F (-479 , 619)
*       1093 = UAC56/F6 (-516 , 639)
*       1093 = UAC58/F (-115.5 , 619)
*       1093 = UAC57/U206/B (-155.5 , 610.5)
*       1093 = UAC57/F6 (-151.5 , 639)
*       1093 = UAC58/U206/B (208 , 610.5)
*       1093 = UAC58/F6 (212 , 639)
*       1101 = UAC55/U218/B (-1007.5 , 566.5)
*       1101 = UAC55/U229/Vout (-968.5 , 568)
*       1102 = UAC55/U222/B (-1014 , 610.5)
*       1102 = UAC55/U206/A (-957 , 615.5)
*       1102 = UAC55/A6 (-955.5 , 645)
*       1102 = UAC52/S (-847 , 689)
*       1102 = UAC52/U218/Vout (-681.5 , 741)
*       1103 = UAC55/U222/Vout (-1052 , 622.5)
*       1103 = UAC55/U218/A (-1081 , 571.5)
*       1111 = UAC55/U262/vout (-1120 , 612.5)
*       1111 = UAC55/U222/A (-1087.5 , 615.5)
*       1112 = UAC55/U238/B (-1143 , 566.5)
*       1112 = UAC55/U220/A (-997.5 , 610.5)
*       1112 = UAC56/U254/Vout (-675 , 524)
*       1112 = UAC56/P (-674 , 497)
*       1112 = UAC55/U236/B (-872 , 566.5)
*       1112 = UAC55/C (-831.5 , 593.5)
*       1112 = UAC55/C6 (-997.5 , 642.5)
*       1113 = UAC55/U245/Vout (-1102.5 , 568)
*       1113 = UAC55/U253/A (-1008.5 , 512.5)
*       1114 = UAC55/U245/Vin (-1116.5 , 568)
*       1114 = UAC55/U238/OUT (-1156 , 555)
*       1115 = UAC55/U262/vin (-1105.5 , 611)
*       1115 = UAC55/U219/OUT (-1155.5 , 599)
*       1121 = UAC85/U229/Vin (-1354 , 568)
*       1121 = UAC85/U220/OUT (-1355.5 , 599)
*       1128 = UAC85/U206/Vout (-1293 , 622.5)
*       1128 = UAC85/U236/A (-1270 , 566.5)
*       1128 = UAC85/U235/B (-1288 , 566.5)
*       1136 = UAC85/U245/Vout (-1474 , 568)
*       1136 = UAC85/U253/A (-1380 , 512.5)
*       1137 = UAC85/U222/Vout (-1423.5 , 622.5)
*       1137 = UAC85/U218/A (-1452.5 , 571.5)
*       1140 = UAC85/U218/B (-1379 , 566.5)
*       1140 = UAC85/U229/Vout (-1340 , 568)
*       1146 = UAC85/U222/B (-1385.5 , 610.5)
*       1146 = UAC85/U206/A (-1328.5 , 615.5)
*       1146 = UAC85/A6 (-1327 , 645)
*       1146 = UAC51/S (-1210.5 , 689)
*       1146 = UAC51/U218/Vout (-1045 , 741)
*       1147 = UAC85/U262/vout (-1491.5 , 612.5)
*       1147 = UAC85/U222/A (-1459 , 615.5)
*       1148 = UAC85/U238/B (-1514.5 , 566.5)
*       1148 = UAC85/U220/A (-1369 , 610.5)
*       1148 = UAC55/U254/Vout (-1038.5 , 524)
*       1148 = UAC55/P (-1037.5 , 497)
*       1148 = UAC85/U236/B (-1243.5 , 566.5)
*       1148 = UAC85/C (-1203 , 593.5)
*       1148 = UAC85/C6 (-1369 , 642.5)
*       1149 = UAC85/U238/OUT (-1527.5 , 555)
*       1149 = UAC85/U245/Vin (-1488 , 568)
*       1150 = UAC85/U219/OUT (-1527 , 599)
*       1150 = UAC85/U262/vin (-1477 , 611)
*       1156 = UAC87/U206/Vout (-1661 , 622.5)
*       1156 = UAC87/U236/A (-1638 , 566.5)
*       1156 = UAC87/U235/B (-1656 , 566.5)
*       1163 = UAC87/U218/B (-1747 , 566.5)
*       1163 = UAC87/U229/Vout (-1708 , 568)
*       1164 = UAC87/U229/Vin (-1722 , 568)
*       1164 = UAC87/U220/OUT (-1723.5 , 599)
*       1165 = UAC87/U222/B (-1753.5 , 610.5)
*       1165 = UAC87/U206/A (-1696.5 , 615.5)
*       1165 = UAC87/A6 (-1695 , 645)
*       1165 = UAC81/S (-1582 , 689)
*       1165 = UAC81/U218/Vout (-1416.5 , 741)
*       1177 = UAC87/U262/vout (-1859.5 , 612.5)
*       1177 = UAC87/U222/A (-1827 , 615.5)
*       1178 = UAC87/U245/Vout (-1842 , 568)
*       1178 = UAC87/U253/A (-1748 , 512.5)
*       1180 = UAC87/U218/A (-1820.5 , 571.5)
*       1180 = UAC87/U222/Vout (-1791.5 , 622.5)
*       1183 = UAC87/U238/OUT (-1895.5 , 555)
*       1183 = UAC87/U245/Vin (-1856 , 568)
*       1184 = UAC87/U219/OUT (-1895 , 599)
*       1184 = UAC87/U262/vin (-1845 , 611)
*       1187 = UAC87/U238/B (-1882.5 , 566.5)
*       1187 = UAC87/U220/A (-1737 , 610.5)
*       1187 = UAC87/U236/B (-1611.5 , 566.5)
*       1187 = UAC85/U254/Vout (-1410 , 524)
*       1187 = UAC85/P (-1409 , 497)
*       1187 = UAC87/C (-1571 , 593.5)
*       1187 = UAC87/C6 (-1737 , 642.5)
*       1191 = UAC88/U206/Vout (-2025 , 622.5)
*       1191 = UAC88/U236/A (-2002 , 566.5)
*       1191 = UAC88/U235/B (-2020 , 566.5)
*       1195 = UAC88/U246/Vin (-1994 , 524)
*       1195 = UAC88/U236/OUT (-1988.5 , 555)
*       1205 = UAC88/U218/B (-2111 , 566.5)
*       1205 = UAC88/U229/Vout (-2072 , 568)
*       1206 = UAC88/U222/B (-2117.5 , 610.5)
*       1206 = UAC88/U206/A (-2060.5 , 615.5)
*       1206 = UAC88/A6 (-2059 , 645)
*       1206 = UAC82/S (-1950.5 , 689)
*       1206 = UAC82/U218/Vout (-1785 , 741)
*       1207 = UAC88/U222/Vout (-2155.5 , 622.5)
*       1207 = UAC88/U218/A (-2184.5 , 571.5)
*       1213 = UAC88/U229/Vin (-2086 , 568)
*       1213 = UAC88/U220/OUT (-2087.5 , 599)
*       1217 = UAC88/U262/vout (-2223.5 , 612.5)
*       1217 = UAC88/U222/A (-2191 , 615.5)
*       1218 = UAC88/U238/B (-2246.5 , 566.5)
*       1218 = UAC88/U220/A (-2101 , 610.5)
*       1218 = UAC87/U254/Vout (-1778 , 524)
*       1218 = UAC87/P (-1777 , 497)
*       1218 = UAC88/U236/B (-1975.5 , 566.5)
*       1218 = UAC88/C (-1935 , 593.5)
*       1218 = UAC88/C6 (-2101 , 642.5)
*       1219 = UAC88/U245/Vout (-2206 , 568)
*       1219 = UAC88/U253/A (-2112 , 512.5)
*       1220 = UAC88/U245/Vin (-2220 , 568)
*       1220 = UAC88/U238/OUT (-2259.5 , 555)
*       1221 = UAC88/U262/vin (-2209 , 611)
*       1221 = UAC88/U219/OUT (-2259 , 599)
*       1227 = UAC90/U229/Vin (-2456.5 , 568)
*       1227 = UAC90/U220/OUT (-2458 , 599)
*       1234 = UAC90/U206/Vout (-2395.5 , 622.5)
*       1234 = UAC90/U236/A (-2372.5 , 566.5)
*       1234 = UAC90/U235/B (-2390.5 , 566.5)
*       1241 = UAC90/U222/B (-2488 , 610.5)
*       1241 = UAC90/U206/A (-2431 , 615.5)
*       1241 = UAC90/A6 (-2429.5 , 645)
*       1241 = UAC84/S (-2314 , 689)
*       1241 = UAC84/U218/Vout (-2148.5 , 741)
*       1244 = UAC90/U245/Vout (-2576.5 , 568)
*       1244 = UAC90/U253/A (-2482.5 , 512.5)
*       1245 = UAC90/U222/Vout (-2526 , 622.5)
*       1245 = UAC90/U218/A (-2555 , 571.5)
*       1247 = UAC90/U218/B (-2481.5 , 566.5)
*       1247 = UAC90/U229/Vout (-2442.5 , 568)
*       1253 = UAC90/U262/vout (-2594 , 612.5)
*       1253 = UAC90/U222/A (-2561.5 , 615.5)
*       1254 = UAC90/U238/B (-2617 , 566.5)
*       1254 = UAC90/U220/A (-2471.5 , 610.5)
*       1254 = UAC88/U254/Vout (-2142 , 524)
*       1254 = UAC88/P (-2141 , 497)
*       1254 = UAC90/U236/B (-2346 , 566.5)
*       1254 = UAC90/C (-2305.5 , 593.5)
*       1254 = UAC90/C6 (-2471.5 , 642.5)
*       1255 = UAC90/U238/OUT (-2630 , 555)
*       1255 = UAC90/U245/Vin (-2590.5 , 568)
*       1256 = UAC90/U219/OUT (-2629.5 , 599)
*       1256 = UAC90/U262/vin (-2579.5 , 611)
*       1259 = UAC118/U229/OUT (-2905.5 , 553.5)
*       1259 = UAC118/U230/vin (-2875 , 565)
*       1260 = UAC118/U228/vin (-2896 , 610.5)
*       1260 = UAC118/U227/O/P (-2911.5 , 618.5)
*       1261 = UAC118/U227/B (-2925 , 625)
*       1261 = UAC118/U226/vout (-2930.5 , 564)
*       1266 = UAC118/U222/OUT (-3018.5 , 599)
*       1266 = UAC118/U223/vin (-2988 , 610.5)
*       1267 = UAC118/U225/A (-3003 , 565)
*       1267 = UAC118/U224/vout (-3014.5 , 564)
*       1269 = UAC118/U222/B (-3005.5 , 610.5)
*       1269 = UAC118/U225/B (-2976.5 , 565)
*       1269 = UAC118/L (-3006.5 , 648)
*       1269 = Lf3 (-3006 , 655)
*       1271 = UAC118/U226/vin (-2959 , 565)
*       1271 = UAC118/U225/OUT (-2989.5 , 553.5)
*       1275 = UAC58/U247/Vin (153 , 524)
*       1275 = UAC58/U235/OUT (162 , 555)
*       1276 = UAC58/U246/Vin (201 , 524)
*       1276 = UAC58/U236/OUT (206.5 , 555)
*       1277 = UAC58/U253/C (123 , 512.5)
*       1277 = UAC58/U247/Vout (167 , 524)
*       1284 = UAC61/U222/B (77 , 448)
*       1284 = UAC119/U223/vout (-3334 , 447)
*       1284 = UAC119/An (-3335 , 491)
*       1284 = UAC61/U206/A (134 , 453)
*       1284 = UAC61/A6 (135.5 , 482.5)
*       1285 = UAC58/U254/Vin (39 , 524)
*       1285 = UAC58/U253/OUT (73.5 , 512.5)
*       1286 = UAC58/U253/B (95.5 , 513)
*       1286 = UAC58/U246/Vout (215 , 524)
*       1287 = UAC119/U228/vout (-3242 , 447)
*       1287 = UAC119/D (-3205.5 , 442.5)
*       1287 = UAC119/Dn (-3243.5 , 489)
*       1287 = UAC95/D (-3048.5 , 444.5)
*       1287 = UAC95/U219/B (-2984 , 448)
*       1287 = UAC95/D6 (-2984.5 , 475)
*       1287 = UAC95/U220/B (-2812.5 , 448)
*       1287 = UAC94/D (-2681.5 , 444.5)
*       1287 = UAC94/U219/B (-2617 , 448)
*       1287 = UAC94/D6 (-2617.5 , 475)
*       1287 = UAC94/U220/B (-2445.5 , 448)
*       1287 = UAC93/D (-2311 , 444.5)
*       1287 = UAC93/U219/B (-2246.5 , 448)
*       1287 = UAC93/D6 (-2247 , 475)
*       1287 = UAC93/U220/B (-2075 , 448)
*       1287 = UAC92/D (-1947 , 444.5)
*       1287 = UAC92/U219/B (-1882.5 , 448)
*       1287 = UAC92/D6 (-1883 , 475)
*       1287 = UAC92/U220/B (-1711 , 448)
*       1287 = UAC91/D (-1579 , 444.5)
*       1287 = UAC91/U219/B (-1514.5 , 448)
*       1287 = UAC91/D6 (-1515 , 475)
*       1287 = UAC91/U220/B (-1343 , 448)
*       1287 = UAC59/D (-1207.5 , 444.5)
*       1287 = UAC59/U219/B (-1143 , 448)
*       1287 = UAC59/D6 (-1143.5 , 475)
*       1287 = UAC59/U220/B (-971.5 , 448)
*       1287 = UAC66/D (-844 , 444.5)
*       1287 = UAC66/U219/B (-779.5 , 448)
*       1287 = UAC66/D6 (-780 , 475)
*       1287 = UAC66/U220/B (-608 , 448)
*       1287 = UAC60/D (-479.5 , 444.5)
*       1287 = UAC60/U219/B (-415 , 448)
*       1287 = UAC60/D6 (-415.5 , 475)
*       1287 = UAC60/U220/B (-243.5 , 448)
*       1287 = UAC61/D (-116 , 444.5)
*       1287 = UAC61/U219/B (-51.5 , 448)
*       1287 = UAC61/D6 (-52 , 475)
*       1287 = UAC61/U220/B (120 , 448)
*       1292 = UAC61/U262/vout (-29 , 450)
*       1292 = UAC61/U222/A (3.5 , 453)
*       1293 = UAC61/U219/OUT (-64.5 , 436.5)
*       1293 = UAC61/U262/vin (-14.5 , 448.5)
*       1295 = UAC60/U206/A (-229.5 , 453)
*       1295 = UAC60/A6 (-228 , 482.5)
*       1295 = UAC60/U222/B (-286.5 , 448)
*       1295 = UAC58/S (-119.5 , 526.5)
*       1295 = UAC58/U218/Vout (46 , 578.5)
*       1296 = UAC57/U246/Vin (-162.5 , 524)
*       1296 = UAC57/U236/OUT (-157 , 555)
*       1299 = UAC57/U253/B (-268 , 513)
*       1299 = UAC57/U246/Vout (-148.5 , 524)
*       1300 = UAC57/U247/Vin (-210.5 , 524)
*       1300 = UAC57/U235/OUT (-201.5 , 555)
*       1301 = UAC57/U253/C (-240.5 , 512.5)
*       1301 = UAC57/U247/Vout (-196.5 , 524)
*       1305 = UAC60/U206/Vout (-194 , 460)
*       1305 = UAC60/U236/A (-171 , 404)
*       1305 = UAC60/U235/B (-189 , 404)
*       1311 = UAC57/U254/Vin (-324.5 , 524)
*       1311 = UAC57/U253/OUT (-290 , 512.5)
*       1315 = UAC60/U219/OUT (-428 , 436.5)
*       1315 = UAC60/U262/vin (-378 , 448.5)
*       1316 = UAC60/U262/vout (-392.5 , 450)
*       1316 = UAC60/U222/A (-360 , 453)
*       1317 = UAC66/U206/A (-594 , 453)
*       1317 = UAC66/A6 (-592.5 , 482.5)
*       1317 = UAC66/U222/B (-651 , 448)
*       1317 = UAC57/S (-483 , 526.5)
*       1317 = UAC57/U218/Vout (-317.5 , 578.5)
*       1322 = UAC56/U247/Vin (-575 , 524)
*       1322 = UAC56/U235/OUT (-566 , 555)
*       1323 = UAC56/U246/Vin (-527 , 524)
*       1323 = UAC56/U236/OUT (-521.5 , 555)
*       1327 = UAC56/U254/Vin (-689 , 524)
*       1327 = UAC56/U253/OUT (-654.5 , 512.5)
*       1328 = UAC56/U253/B (-632.5 , 513)
*       1328 = UAC56/U246/Vout (-513 , 524)
*       1329 = UAC56/U253/C (-605 , 512.5)
*       1329 = UAC56/U247/Vout (-561 , 524)
*       1335 = UAC66/U262/vout (-757 , 450)
*       1335 = UAC66/U222/A (-724.5 , 453)
*       1338 = UAC66/U219/OUT (-792.5 , 436.5)
*       1338 = UAC66/U262/vin (-742.5 , 448.5)
*       1339 = UAC59/U222/B (-1014.5 , 448)
*       1339 = UAC59/U206/A (-957.5 , 453)
*       1339 = UAC59/A6 (-956 , 482.5)
*       1339 = UAC56/S (-847.5 , 526.5)
*       1339 = UAC56/U218/Vout (-682 , 578.5)
*       1344 = UAC55/U247/Vin (-938.5 , 524)
*       1344 = UAC55/U235/OUT (-929.5 , 555)
*       1345 = UAC55/U246/Vin (-890.5 , 524)
*       1345 = UAC55/U236/OUT (-885 , 555)
*       1346 = UAC55/U253/C (-968.5 , 512.5)
*       1346 = UAC55/U247/Vout (-924.5 , 524)
*       1349 = UAC119/U220/B (-3241 , 357.5)
*       1349 = UAC119/U230/vout (-3221 , 401.5)
*       1349 = UAC119/Fn (-3205 , 425.5)
*       1349 = UAC95/F (-3048.5 , 456.5)
*       1349 = UAC95/U206/B (-2725 , 448)
*       1349 = UAC95/F6 (-2721 , 476.5)
*       1349 = UAC94/F (-2681.5 , 456.5)
*       1349 = UAC94/U206/B (-2358 , 448)
*       1349 = UAC94/F6 (-2354 , 476.5)
*       1349 = UAC93/F (-2311 , 456.5)
*       1349 = UAC93/U206/B (-1987.5 , 448)
*       1349 = UAC93/F6 (-1983.5 , 476.5)
*       1349 = UAC92/F (-1947 , 456.5)
*       1349 = UAC92/U206/B (-1623.5 , 448)
*       1349 = UAC92/F6 (-1619.5 , 476.5)
*       1349 = UAC91/F (-1579 , 456.5)
*       1349 = UAC91/U206/B (-1255.5 , 448)
*       1349 = UAC91/F6 (-1251.5 , 476.5)
*       1349 = UAC59/F (-1207.5 , 456.5)
*       1349 = UAC66/F (-844 , 456.5)
*       1349 = UAC59/U206/B (-884 , 448)
*       1349 = UAC59/F6 (-880 , 476.5)
*       1349 = UAC66/U206/B (-520.5 , 448)
*       1349 = UAC66/F6 (-516.5 , 476.5)
*       1349 = UAC60/F (-479.5 , 456.5)
*       1349 = UAC61/F (-116 , 456.5)
*       1349 = UAC60/U206/B (-156 , 448)
*       1349 = UAC60/F6 (-152 , 476.5)
*       1349 = UAC61/U206/B (207.5 , 448)
*       1349 = UAC61/F6 (211.5 , 476.5)
*       1355 = UAC55/U254/Vin (-1052.5 , 524)
*       1355 = UAC55/U253/OUT (-1018 , 512.5)
*       1356 = UAC55/U253/B (-996 , 513)
*       1356 = UAC55/U246/Vout (-876.5 , 524)
*       1360 = UAC59/U219/OUT (-1156 , 436.5)
*       1360 = UAC59/U262/vin (-1106 , 448.5)
*       1361 = UAC59/U262/vout (-1120.5 , 450)
*       1361 = UAC59/U222/A (-1088 , 453)
*       1363 = UAC91/U206/A (-1329 , 453)
*       1363 = UAC91/A6 (-1327.5 , 482.5)
*       1363 = UAC91/U222/B (-1386 , 448)
*       1363 = UAC55/S (-1211 , 526.5)
*       1363 = UAC55/U218/Vout (-1045.5 , 578.5)
*       1364 = UAC85/U246/Vin (-1262 , 524)
*       1364 = UAC85/U236/OUT (-1256.5 , 555)
*       1367 = UAC85/U253/B (-1367.5 , 513)
*       1367 = UAC85/U246/Vout (-1248 , 524)
*       1368 = UAC85/U247/Vin (-1310 , 524)
*       1368 = UAC85/U235/OUT (-1301 , 555)
*       1369 = UAC85/U253/C (-1340 , 512.5)
*       1369 = UAC85/U247/Vout (-1296 , 524)
*       1373 = UAC91/U206/Vout (-1293.5 , 460)
*       1373 = UAC91/U236/A (-1270.5 , 404)
*       1373 = UAC91/U235/B (-1288.5 , 404)
*       1379 = UAC85/U254/Vin (-1424 , 524)
*       1379 = UAC85/U253/OUT (-1389.5 , 512.5)
*       1383 = UAC91/U219/OUT (-1527.5 , 436.5)
*       1383 = UAC91/U262/vin (-1477.5 , 448.5)
*       1384 = UAC91/U262/vout (-1492 , 450)
*       1384 = UAC91/U222/A (-1459.5 , 453)
*       1385 = UAC92/U206/A (-1697 , 453)
*       1385 = UAC92/A6 (-1695.5 , 482.5)
*       1385 = UAC92/U222/B (-1754 , 448)
*       1385 = UAC85/S (-1582.5 , 526.5)
*       1385 = UAC85/U218/Vout (-1417 , 578.5)
*       1390 = UAC87/U247/Vin (-1678 , 524)
*       1390 = UAC87/U235/OUT (-1669 , 555)
*       1391 = UAC87/U246/Vin (-1630 , 524)
*       1391 = UAC87/U236/OUT (-1624.5 , 555)
*       1395 = UAC87/U253/B (-1735.5 , 513)
*       1395 = UAC87/U246/Vout (-1616 , 524)
*       1396 = UAC87/U253/C (-1708 , 512.5)
*       1396 = UAC87/U247/Vout (-1664 , 524)
*       1401 = UAC92/U262/vout (-1860 , 450)
*       1401 = UAC92/U222/A (-1827.5 , 453)
*       1402 = UAC87/U254/Vin (-1792 , 524)
*       1402 = UAC87/U253/OUT (-1757.5 , 512.5)
*       1404 = UAC92/U218/A (-1821 , 409)
*       1404 = UAC92/U222/Vout (-1792 , 460)
*       1407 = UAC92/U219/OUT (-1895.5 , 436.5)
*       1407 = UAC92/U262/vin (-1845.5 , 448.5)
*       1408 = UAC93/U222/B (-2118 , 448)
*       1408 = UAC93/U206/A (-2061 , 453)
*       1408 = UAC93/A6 (-2059.5 , 482.5)
*       1408 = UAC87/S (-1950.5 , 526.5)
*       1408 = UAC87/U218/Vout (-1785 , 578.5)
*       1413 = UAC88/U247/Vin (-2042 , 524)
*       1413 = UAC88/U235/OUT (-2033 , 555)
*       1414 = UAC88/U253/C (-2072 , 512.5)
*       1414 = UAC88/U247/Vout (-2028 , 524)
*       1421 = UAC88/U254/Vin (-2156 , 524)
*       1421 = UAC88/U253/OUT (-2121.5 , 512.5)
*       1422 = UAC88/U253/B (-2099.5 , 513)
*       1422 = UAC88/U246/Vout (-1980 , 524)
*       1425 = UAC93/U229/Vin (-2086.5 , 405.5)
*       1425 = UAC93/U220/OUT (-2088 , 436.5)
*       1428 = UAC93/U219/OUT (-2259.5 , 436.5)
*       1428 = UAC93/U262/vin (-2209.5 , 448.5)
*       1429 = UAC93/U262/vout (-2224 , 450)
*       1429 = UAC93/U222/A (-2191.5 , 453)
*       1431 = UAC94/U206/A (-2431.5 , 453)
*       1431 = UAC94/A6 (-2430 , 482.5)
*       1431 = UAC94/U222/B (-2488.5 , 448)
*       1431 = UAC88/S (-2314.5 , 526.5)
*       1431 = UAC88/U218/Vout (-2149 , 578.5)
*       1432 = UAC90/U246/Vin (-2364.5 , 524)
*       1432 = UAC90/U236/OUT (-2359 , 555)
*       1435 = UAC90/U253/B (-2470 , 513)
*       1435 = UAC90/U246/Vout (-2350.5 , 524)
*       1436 = UAC90/U247/Vin (-2412.5 , 524)
*       1436 = UAC90/U235/OUT (-2403.5 , 555)
*       1437 = UAC90/U253/C (-2442.5 , 512.5)
*       1437 = UAC90/U247/Vout (-2398.5 , 524)
*       1441 = UAC94/U206/Vout (-2396 , 460)
*       1441 = UAC94/U236/A (-2373 , 404)
*       1441 = UAC94/U235/B (-2391 , 404)
*       1447 = UAC90/U254/Vin (-2526.5 , 524)
*       1447 = UAC90/U253/OUT (-2492 , 512.5)
*       1451 = UAC94/U262/vout (-2594.5 , 450)
*       1451 = UAC94/U222/A (-2562 , 453)
*       1452 = UAC95/U206/A (-2798.5 , 453)
*       1452 = UAC95/A6 (-2797 , 482.5)
*       1452 = UAC95/U222/B (-2855.5 , 448)
*       1452 = UAC90/S (-2685 , 526.5)
*       1452 = UAC90/U218/Vout (-2519.5 , 578.5)
*       1454 = UAC94/U219/OUT (-2630 , 436.5)
*       1454 = UAC94/U262/vin (-2580 , 448.5)
*       1465 = UAC95/U262/vout (-2961.5 , 450)
*       1465 = UAC95/U222/A (-2929 , 453)
*       1469 = UAC118/U220/A (-2940 , 525)
*       1469 = UAC118/U232/vout (-2951.5 , 519)
*       1472 = UAC95/U218/A (-2922.5 , 409)
*       1472 = UAC95/U222/Vout (-2893.5 , 460)
*       1475 = UAC118/U231/B (-2997.5 , 520)
*       1475 = UAC118/Pn (-2998 , 493.5)
*       1475 = UAC90/U254/Vout (-2512.5 , 524)
*       1475 = UAC90/P (-2511.5 , 497)
*       1476 = UAC118/U231/OUT (-3010.5 , 508.5)
*       1476 = UAC118/U232/vin (-2980 , 520)
*       1477 = UAC95/U219/OUT (-2997 , 436.5)
*       1477 = UAC95/U262/vin (-2947 , 448.5)
*       1480 = UAC119/U228/vin (-3270.5 , 448)
*       1480 = UAC119/U227/O/P (-3286 , 456)
*       1481 = Q3 (-3312.5 , 523.5)
*       1481 = UAC119/Fn (-3445 , 414)
*       1481 = UAC119/U229/B (-3267 , 402.5)
*       1481 = UAC119/F (-3263.5 , 488)
*       1481 = UAC118/Qn (-3070 , 523)
*       1481 = UAC118/U220/Vout (-2904.5 , 532)
*       1483 = UAC119/U222/OUT (-3393 , 436.5)
*       1483 = UAC119/U223/vin (-3362.5 , 448)
*       1484 = UAC119/U225/B (-3351 , 402.5)
*       1484 = UAC119/U222/B (-3380 , 448)
*       1484 = UAC119/L (-3381 , 485.5)
*       1484 = Lf2 (-3380 , 491)
*       1486 = UAC61/U253/C (122.5 , 350)
*       1486 = UAC61/U247/Vout (166.5 , 361.5)
*       1487 = UAC61/U247/Vin (152.5 , 361.5)
*       1487 = UAC61/U235/OUT (161.5 , 392.5)
*       1488 = UAC61/U246/Vin (200.5 , 361.5)
*       1488 = UAC61/U236/OUT (206 , 392.5)
*       1489 = UAC61/U236/A (192.5 , 404)
*       1489 = UAC61/U235/B (174.5 , 404)
*       1489 = UAC61/U206/Vout (169.5 , 460)
*       1495 = UAC61/U218/B (83.5 , 404)
*       1495 = UAC61/U229/Vout (122.5 , 405.5)
*       1496 = UAC61/U254/Vin (38.5 , 361.5)
*       1496 = UAC61/U253/OUT (73 , 350)
*       1497 = UAC61/U253/B (95 , 350.5)
*       1497 = UAC61/U246/Vout (214.5 , 361.5)
*       1498 = UAC61/U229/Vin (108.5 , 405.5)
*       1498 = UAC61/U220/OUT (107 , 436.5)
*       1499 = UAC61/U218/A (10 , 409)
*       1499 = UAC61/U222/Vout (39 , 460)
*       1505 = UAC61/U245/Vout (-11.5 , 405.5)
*       1505 = UAC61/U253/A (82.5 , 350)
*       1506 = UAC61/U245/Vin (-25.5 , 405.5)
*       1506 = UAC61/U238/OUT (-65 , 392.5)
*       1508 = UAC60/U246/Vin (-163 , 361.5)
*       1508 = UAC60/U236/OUT (-157.5 , 392.5)
*       1510 = UAC60/U253/B (-268.5 , 350.5)
*       1510 = UAC60/U246/Vout (-149 , 361.5)
*       1511 = UAC60/U253/C (-241 , 350)
*       1511 = UAC60/U247/Vout (-197 , 361.5)
*       1512 = UAC60/U247/Vin (-211 , 361.5)
*       1512 = UAC60/U235/OUT (-202 , 392.5)
*       1513 = UAC60/U229/Vin (-255 , 405.5)
*       1513 = UAC60/U220/OUT (-256.5 , 436.5)
*       1520 = UAC60/U245/Vout (-375 , 405.5)
*       1520 = UAC60/U253/A (-281 , 350)
*       1521 = UAC60/U254/Vin (-325 , 361.5)
*       1521 = UAC60/U253/OUT (-290.5 , 350)
*       1522 = UAC60/U218/A (-353.5 , 409)
*       1522 = UAC60/U222/Vout (-324.5 , 460)
*       1524 = UAC60/U218/B (-280 , 404)
*       1524 = UAC60/U229/Vout (-241 , 405.5)
*       1527 = UAC60/U238/OUT (-428.5 , 392.5)
*       1527 = UAC60/U245/Vin (-389 , 405.5)
*       1528 = UAC60/U238/B (-415.5 , 404)
*       1528 = UAC60/U220/A (-270 , 448)
*       1528 = UAC60/C6 (-270 , 480)
*       1528 = UAC61/U254/Vout (52.5 , 361.5)
*       1528 = UAC61/P (53.5 , 334.5)
*       1528 = UAC60/U236/B (-144.5 , 404)
*       1528 = UAC60/C (-104 , 431)
*       1530 = UAC66/U247/Vin (-575.5 , 361.5)
*       1530 = UAC66/U235/OUT (-566.5 , 392.5)
*       1531 = UAC66/U246/Vin (-527.5 , 361.5)
*       1531 = UAC66/U236/OUT (-522 , 392.5)
*       1532 = UAC66/U236/A (-535.5 , 404)
*       1532 = UAC66/U235/B (-553.5 , 404)
*       1532 = UAC66/U206/Vout (-558.5 , 460)
*       1536 = UAC66/U218/B (-644.5 , 404)
*       1536 = UAC66/U229/Vout (-605.5 , 405.5)
*       1537 = UAC66/U253/B (-633 , 350.5)
*       1537 = UAC66/U246/Vout (-513.5 , 361.5)
*       1538 = UAC66/U253/C (-605.5 , 350)
*       1538 = UAC66/U247/Vout (-561.5 , 361.5)
*       1539 = UAC66/U229/Vin (-619.5 , 405.5)
*       1539 = UAC66/U220/OUT (-621 , 436.5)
*       1547 = UAC66/U245/Vout (-739.5 , 405.5)
*       1547 = UAC66/U253/A (-645.5 , 350)
*       1548 = UAC66/U254/Vin (-689.5 , 361.5)
*       1548 = UAC66/U253/OUT (-655 , 350)
*       1549 = UAC66/U218/A (-718 , 409)
*       1549 = UAC66/U222/Vout (-689 , 460)
*       1550 = UAC66/U238/OUT (-793 , 392.5)
*       1550 = UAC66/U245/Vin (-753.5 , 405.5)
*       1552 = UAC66/U238/B (-780 , 404)
*       1552 = UAC66/U220/A (-634.5 , 448)
*       1552 = UAC66/C6 (-634.5 , 480)
*       1552 = UAC66/U236/B (-509 , 404)
*       1552 = UAC60/U254/Vout (-311 , 361.5)
*       1552 = UAC60/P (-310 , 334.5)
*       1552 = UAC66/C (-468.5 , 431)
*       1554 = UAC59/U253/C (-969 , 350)
*       1554 = UAC59/U247/Vout (-925 , 361.5)
*       1555 = UAC59/U247/Vin (-939 , 361.5)
*       1555 = UAC59/U235/OUT (-930 , 392.5)
*       1556 = UAC59/U246/Vin (-891 , 361.5)
*       1556 = UAC59/U236/OUT (-885.5 , 392.5)
*       1557 = UAC59/U236/A (-899 , 404)
*       1557 = UAC59/U235/B (-917 , 404)
*       1557 = UAC59/U206/Vout (-922 , 460)
*       1558 = UAC59/U229/Vin (-983 , 405.5)
*       1558 = UAC59/U220/OUT (-984.5 , 436.5)
*       1564 = UAC59/U218/B (-1008 , 404)
*       1564 = UAC59/U229/Vout (-969 , 405.5)
*       1565 = UAC59/U254/Vin (-1053 , 361.5)
*       1565 = UAC59/U253/OUT (-1018.5 , 350)
*       1566 = UAC59/U218/A (-1081.5 , 409)
*       1566 = UAC59/U222/Vout (-1052.5 , 460)
*       1568 = UAC59/U253/B (-996.5 , 350.5)
*       1568 = UAC59/U246/Vout (-877 , 361.5)
*       1572 = UAC59/U245/Vout (-1103 , 405.5)
*       1572 = UAC59/U253/A (-1009 , 350)
*       1573 = UAC59/U245/Vin (-1117 , 405.5)
*       1573 = UAC59/U238/OUT (-1156.5 , 392.5)
*       1574 = UAC59/U238/B (-1143.5 , 404)
*       1574 = UAC59/U220/A (-998 , 448)
*       1574 = UAC59/C6 (-998 , 480)
*       1574 = UAC66/U254/Vout (-675.5 , 361.5)
*       1574 = UAC66/P (-674.5 , 334.5)
*       1574 = UAC59/U236/B (-872.5 , 404)
*       1574 = UAC59/C (-832 , 431)
*       1576 = UAC91/U246/Vin (-1262.5 , 361.5)
*       1576 = UAC91/U236/OUT (-1257 , 392.5)
*       1578 = UAC91/U253/B (-1368 , 350.5)
*       1578 = UAC91/U246/Vout (-1248.5 , 361.5)
*       1579 = UAC91/U253/C (-1340.5 , 350)
*       1579 = UAC91/U247/Vout (-1296.5 , 361.5)
*       1580 = UAC91/U247/Vin (-1310.5 , 361.5)
*       1580 = UAC91/U235/OUT (-1301.5 , 392.5)
*       1581 = UAC91/U229/Vin (-1354.5 , 405.5)
*       1581 = UAC91/U220/OUT (-1356 , 436.5)
*       1588 = UAC91/U245/Vout (-1474.5 , 405.5)
*       1588 = UAC91/U253/A (-1380.5 , 350)
*       1589 = UAC91/U254/Vin (-1424.5 , 361.5)
*       1589 = UAC91/U253/OUT (-1390 , 350)
*       1590 = UAC91/U218/A (-1453 , 409)
*       1590 = UAC91/U222/Vout (-1424 , 460)
*       1592 = UAC91/U218/B (-1379.5 , 404)
*       1592 = UAC91/U229/Vout (-1340.5 , 405.5)
*       1595 = UAC91/U238/OUT (-1528 , 392.5)
*       1595 = UAC91/U245/Vin (-1488.5 , 405.5)
*       1596 = UAC91/U238/B (-1515 , 404)
*       1596 = UAC91/U220/A (-1369.5 , 448)
*       1596 = UAC91/C6 (-1369.5 , 480)
*       1596 = UAC59/U254/Vout (-1039 , 361.5)
*       1596 = UAC59/P (-1038 , 334.5)
*       1596 = UAC91/U236/B (-1244 , 404)
*       1596 = UAC91/C (-1203.5 , 431)
*       1598 = UAC92/U247/Vin (-1678.5 , 361.5)
*       1598 = UAC92/U235/OUT (-1669.5 , 392.5)
*       1599 = UAC92/U246/Vin (-1630.5 , 361.5)
*       1599 = UAC92/U236/OUT (-1625 , 392.5)
*       1600 = UAC92/U236/A (-1638.5 , 404)
*       1600 = UAC92/U235/B (-1656.5 , 404)
*       1600 = UAC92/U206/Vout (-1661.5 , 460)
*       1604 = UAC92/U218/B (-1747.5 , 404)
*       1604 = UAC92/U229/Vout (-1708.5 , 405.5)
*       1605 = UAC92/U253/B (-1736 , 350.5)
*       1605 = UAC92/U246/Vout (-1616.5 , 361.5)
*       1606 = UAC92/U253/C (-1708.5 , 350)
*       1606 = UAC92/U247/Vout (-1664.5 , 361.5)
*       1607 = UAC92/U229/Vin (-1722.5 , 405.5)
*       1607 = UAC92/U220/OUT (-1724 , 436.5)
*       1614 = UAC92/U245/Vout (-1842.5 , 405.5)
*       1614 = UAC92/U253/A (-1748.5 , 350)
*       1615 = UAC92/U254/Vin (-1792.5 , 361.5)
*       1615 = UAC92/U253/OUT (-1758 , 350)
*       1617 = UAC92/U238/OUT (-1896 , 392.5)
*       1617 = UAC92/U245/Vin (-1856.5 , 405.5)
*       1619 = UAC92/U238/B (-1883 , 404)
*       1619 = UAC92/U220/A (-1737.5 , 448)
*       1619 = UAC92/C6 (-1737.5 , 480)
*       1619 = UAC92/U236/B (-1612 , 404)
*       1619 = UAC91/U254/Vout (-1410.5 , 361.5)
*       1619 = UAC91/P (-1409.5 , 334.5)
*       1619 = UAC92/C (-1571.5 , 431)
*       1620 = UAC93/U253/C (-2072.5 , 350)
*       1620 = UAC93/U247/Vout (-2028.5 , 361.5)
*       1621 = UAC93/U247/Vin (-2042.5 , 361.5)
*       1621 = UAC93/U235/OUT (-2033.5 , 392.5)
*       1622 = UAC93/U236/A (-2002.5 , 404)
*       1622 = UAC93/U235/B (-2020.5 , 404)
*       1622 = UAC93/U206/Vout (-2025.5 , 460)
*       1625 = UAC93/U246/Vin (-1994.5 , 361.5)
*       1625 = UAC93/U236/OUT (-1989 , 392.5)
*       1629 = UAC93/U218/B (-2111.5 , 404)
*       1629 = UAC93/U229/Vout (-2072.5 , 405.5)
*       1630 = UAC93/U254/Vin (-2156.5 , 361.5)
*       1630 = UAC93/U253/OUT (-2122 , 350)
*       1631 = UAC93/U253/B (-2100 , 350.5)
*       1631 = UAC93/U246/Vout (-1980.5 , 361.5)
*       1632 = UAC93/U218/A (-2185 , 409)
*       1632 = UAC93/U222/Vout (-2156 , 460)
*       1638 = UAC93/U245/Vout (-2206.5 , 405.5)
*       1638 = UAC93/U253/A (-2112.5 , 350)
*       1639 = UAC93/U245/Vin (-2220.5 , 405.5)
*       1639 = UAC93/U238/OUT (-2260 , 392.5)
*       1640 = UAC93/U238/B (-2247 , 404)
*       1640 = UAC93/U220/A (-2101.5 , 448)
*       1640 = UAC93/C6 (-2101.5 , 480)
*       1640 = UAC92/U254/Vout (-1778.5 , 361.5)
*       1640 = UAC92/P (-1777.5 , 334.5)
*       1640 = UAC93/U236/B (-1976 , 404)
*       1640 = UAC93/C (-1935.5 , 431)
*       1642 = UAC94/U246/Vin (-2365 , 361.5)
*       1642 = UAC94/U236/OUT (-2359.5 , 392.5)
*       1644 = UAC94/U253/B (-2470.5 , 350.5)
*       1644 = UAC94/U246/Vout (-2351 , 361.5)
*       1645 = UAC94/U253/C (-2443 , 350)
*       1645 = UAC94/U247/Vout (-2399 , 361.5)
*       1646 = UAC94/U247/Vin (-2413 , 361.5)
*       1646 = UAC94/U235/OUT (-2404 , 392.5)
*       1647 = UAC94/U229/Vin (-2457 , 405.5)
*       1647 = UAC94/U220/OUT (-2458.5 , 436.5)
*       1654 = UAC94/U245/Vout (-2577 , 405.5)
*       1654 = UAC94/U253/A (-2483 , 350)
*       1655 = UAC94/U254/Vin (-2527 , 361.5)
*       1655 = UAC94/U253/OUT (-2492.5 , 350)
*       1656 = UAC94/U218/A (-2555.5 , 409)
*       1656 = UAC94/U222/Vout (-2526.5 , 460)
*       1658 = UAC94/U218/B (-2482 , 404)
*       1658 = UAC94/U229/Vout (-2443 , 405.5)
*       1661 = UAC94/U238/OUT (-2630.5 , 392.5)
*       1661 = UAC94/U245/Vin (-2591 , 405.5)
*       1662 = UAC94/U238/B (-2617.5 , 404)
*       1662 = UAC94/U220/A (-2472 , 448)
*       1662 = UAC94/C6 (-2472 , 480)
*       1662 = UAC93/U254/Vout (-2142.5 , 361.5)
*       1662 = UAC93/P (-2141.5 , 334.5)
*       1662 = UAC94/U236/B (-2346.5 , 404)
*       1662 = UAC94/C (-2306 , 431)
*       1664 = UAC95/U247/Vin (-2780 , 361.5)
*       1664 = UAC95/U235/OUT (-2771 , 392.5)
*       1665 = UAC95/U246/Vin (-2732 , 361.5)
*       1665 = UAC95/U236/OUT (-2726.5 , 392.5)
*       1666 = UAC95/U236/A (-2740 , 404)
*       1666 = UAC95/U235/B (-2758 , 404)
*       1666 = UAC95/U206/Vout (-2763 , 460)
*       1670 = UAC95/U218/B (-2849 , 404)
*       1670 = UAC95/U229/Vout (-2810 , 405.5)
*       1671 = UAC95/U253/B (-2837.5 , 350.5)
*       1671 = UAC95/U246/Vout (-2718 , 361.5)
*       1672 = UAC95/U253/C (-2810 , 350)
*       1672 = UAC95/U247/Vout (-2766 , 361.5)
*       1673 = UAC95/U229/Vin (-2824 , 405.5)
*       1673 = UAC95/U220/OUT (-2825.5 , 436.5)
*       1680 = UAC95/U245/Vout (-2944 , 405.5)
*       1680 = UAC95/U253/A (-2850 , 350)
*       1681 = UAC95/U254/Vin (-2894 , 361.5)
*       1681 = UAC95/U253/OUT (-2859.5 , 350)
*       1683 = UAC95/U238/B (-2984.5 , 404)
*       1683 = UAC95/U220/A (-2839 , 448)
*       1683 = UAC95/C6 (-2839 , 480)
*       1683 = UAC95/U236/B (-2713.5 , 404)
*       1683 = UAC94/U254/Vout (-2513 , 361.5)
*       1683 = UAC94/P (-2512 , 334.5)
*       1683 = UAC95/C (-2673 , 431)
*       1684 = UAC95/U238/OUT (-2997.5 , 392.5)
*       1684 = UAC95/U245/Vin (-2958 , 405.5)
*       1687 = UAC119/U230/vin (-3249.5 , 402.5)
*       1687 = UAC119/U229/OUT (-3280 , 391)
*       1694 = UAC119/U231/B (-3372 , 357.5)
*       1694 = UAC119/Pn (-3372.5 , 331)
*       1694 = UAC95/U254/Vout (-2880 , 361.5)
*       1694 = UAC95/P (-2879 , 334.5)
*       1695 = UAC119/U232/vin (-3354.5 , 357.5)
*       1695 = UAC119/U231/OUT (-3385 , 346)
*       1696 = UAC119/U226/vin (-3333.5 , 402.5)
*       1696 = UAC119/U225/OUT (-3364 , 391)
*       1697 = UAC119/U220/A (-3314.5 , 362.5)
*       1697 = UAC119/U232/vout (-3326 , 356.5)
*       1698 = UAC119/U226/vout (-3305 , 401.5)
*       1698 = UAC119/U227/B (-3299.5 , 462.5)
*       1701 = UAC119/U225/A (-3377.5 , 402.5)
*       1701 = UAC119/U224/vout (-3389 , 401.5)
*       1705 = UAC65/U206/Vout (169 , 297.5)
*       1705 = UAC65/U236/A (192 , 241.5)
*       1705 = UAC65/U235/B (174 , 241.5)
*       1717 = UAC65/U222/B (76.5 , 285.5)
*       1717 = UAC120/U223/vout (-3699 , 284.5)
*       1717 = UAC120/An (-3578.5 , 299)
*       1717 = UAC65/U206/A (133.5 , 290.5)
*       1717 = UAC65/A6 (135 , 320)
*       1718 = UAC65/U229/Vin (108 , 243)
*       1718 = UAC65/U220/OUT (106.5 , 274)
*       1719 = UAC65/U222/Vout (38.5 , 297.5)
*       1719 = UAC65/U218/A (9.5 , 246.5)
*       1721 = UAC120/U228/vout (-3607 , 284.5)
*       1721 = UAC120/D (-3570.5 , 280)
*       1721 = UAC101/D (-3420.5 , 282)
*       1721 = UAC101/U219/B (-3356 , 285.5)
*       1721 = UAC101/D6 (-3356.5 , 312.5)
*       1721 = UAC101/U220/B (-3184.5 , 285.5)
*       1721 = UAC100/D (-3049 , 282)
*       1721 = UAC100/U219/B (-2984.5 , 285.5)
*       1721 = UAC100/D6 (-2985 , 312.5)
*       1721 = UAC100/U220/B (-2813 , 285.5)
*       1721 = UAC99/D (-2682 , 282)
*       1721 = UAC99/U219/B (-2617.5 , 285.5)
*       1721 = UAC99/D6 (-2618 , 312.5)
*       1721 = UAC99/U220/B (-2446 , 285.5)
*       1721 = UAC98/D (-2311.5 , 282)
*       1721 = UAC98/U219/B (-2247 , 285.5)
*       1721 = UAC98/D6 (-2247.5 , 312.5)
*       1721 = UAC98/U220/B (-2075.5 , 285.5)
*       1721 = UAC97/D (-1947.5 , 282)
*       1721 = UAC97/U219/B (-1883 , 285.5)
*       1721 = UAC97/D6 (-1883.5 , 312.5)
*       1721 = UAC97/U220/B (-1711.5 , 285.5)
*       1721 = UAC96/D (-1579.5 , 282)
*       1721 = UAC96/U219/B (-1515 , 285.5)
*       1721 = UAC96/D6 (-1515.5 , 312.5)
*       1721 = UAC96/U220/B (-1343.5 , 285.5)
*       1721 = UAC62/D (-1208 , 282)
*       1721 = UAC62/U219/B (-1143.5 , 285.5)
*       1721 = UAC62/D6 (-1144 , 312.5)
*       1721 = UAC62/U220/B (-972 , 285.5)
*       1721 = UAC63/D (-844.5 , 282)
*       1721 = UAC63/U219/B (-780 , 285.5)
*       1721 = UAC63/D6 (-780.5 , 312.5)
*       1721 = UAC63/U220/B (-608.5 , 285.5)
*       1721 = UAC64/D (-480 , 282)
*       1721 = UAC64/U219/B (-415.5 , 285.5)
*       1721 = UAC64/D6 (-416 , 312.5)
*       1721 = UAC64/U220/B (-244 , 285.5)
*       1721 = UAC65/D (-116.5 , 282)
*       1721 = UAC65/U219/B (-52 , 285.5)
*       1721 = UAC65/D6 (-52.5 , 312.5)
*       1721 = UAC65/U220/B (119.5 , 285.5)
*       1721 = UAC120/Dn (-3608.5 , 326.5)
*       1728 = UAC65/U262/vout (-29.5 , 287.5)
*       1728 = UAC65/U222/A (3 , 290.5)
*       1729 = UAC65/U219/OUT (-65 , 274)
*       1729 = UAC65/U262/vin (-15 , 286)
*       1730 = UAC65/U245/Vout (-12 , 243)
*       1730 = UAC65/U253/A (82 , 187.5)
*       1736 = UAC64/U229/Vin (-255.5 , 243)
*       1736 = UAC64/U220/OUT (-257 , 274)
*       1741 = UAC64/U206/Vout (-194.5 , 297.5)
*       1741 = UAC64/U236/A (-171.5 , 241.5)
*       1741 = UAC64/U235/B (-189.5 , 241.5)
*       1747 = UAC64/U206/A (-230 , 290.5)
*       1747 = UAC64/A6 (-228.5 , 320)
*       1747 = UAC64/U222/B (-287 , 285.5)
*       1747 = UAC61/S (-120 , 364)
*       1747 = UAC61/U218/Vout (45.5 , 416)
*       1751 = UAC64/U222/Vout (-325 , 297.5)
*       1751 = UAC64/U218/A (-354 , 246.5)
*       1753 = UAC64/U218/B (-280.5 , 241.5)
*       1753 = UAC64/U229/Vout (-241.5 , 243)
*       1759 = UAC64/U219/OUT (-428.5 , 274)
*       1759 = UAC64/U262/vin (-378.5 , 286)
*       1760 = UAC64/U262/vout (-393 , 287.5)
*       1760 = UAC64/U222/A (-360.5 , 290.5)
*       1761 = UAC64/U238/B (-416 , 241.5)
*       1761 = UAC64/U220/A (-270.5 , 285.5)
*       1761 = UAC64/C6 (-270.5 , 317.5)
*       1761 = UAC65/U254/Vout (52 , 199)
*       1761 = UAC65/P (53 , 172)
*       1761 = UAC64/U236/B (-145 , 241.5)
*       1761 = UAC64/C (-104.5 , 268.5)
*       1767 = UAC63/U206/Vout (-559 , 297.5)
*       1767 = UAC63/U236/A (-536 , 241.5)
*       1767 = UAC63/U235/B (-554 , 241.5)
*       1774 = UAC63/U206/A (-594.5 , 290.5)
*       1774 = UAC63/A6 (-593 , 320)
*       1774 = UAC63/U222/B (-651.5 , 285.5)
*       1774 = UAC60/S (-483.5 , 364)
*       1774 = UAC60/U218/Vout (-318 , 416)
*       1775 = UAC63/U229/Vin (-620 , 243)
*       1775 = UAC63/U220/OUT (-621.5 , 274)
*       1786 = UAC63/U262/vout (-757.5 , 287.5)
*       1786 = UAC63/U222/A (-725 , 290.5)
*       1787 = UAC63/U218/A (-718.5 , 246.5)
*       1787 = UAC63/U222/Vout (-689.5 , 297.5)
*       1790 = UAC63/U219/OUT (-793 , 274)
*       1790 = UAC63/U262/vin (-743 , 286)
*       1793 = UAC63/U238/B (-780.5 , 241.5)
*       1793 = UAC63/U220/A (-635 , 285.5)
*       1793 = UAC63/C6 (-635 , 317.5)
*       1793 = UAC63/U236/B (-509.5 , 241.5)
*       1793 = UAC64/U254/Vout (-311.5 , 199)
*       1793 = UAC64/P (-310.5 , 172)
*       1793 = UAC63/C (-469 , 268.5)
*       1798 = UAC62/U206/Vout (-922.5 , 297.5)
*       1798 = UAC62/U236/A (-899.5 , 241.5)
*       1798 = UAC62/U235/B (-917.5 , 241.5)
*       1799 = UAC62/U229/Vin (-983.5 , 243)
*       1799 = UAC62/U220/OUT (-985 , 274)
*       1805 = UAC120/U220/B (-3606 , 195)
*       1805 = UAC120/U230/vout (-3586 , 239)
*       1805 = UAC120/Fn (-3570 , 263)
*       1805 = UAC101/F (-3420.5 , 294)
*       1805 = UAC101/U206/B (-3097 , 285.5)
*       1805 = UAC101/F6 (-3093 , 314)
*       1805 = UAC100/F (-3049 , 294)
*       1805 = UAC100/U206/B (-2725.5 , 285.5)
*       1805 = UAC100/F6 (-2721.5 , 314)
*       1805 = UAC99/F (-2682 , 294)
*       1805 = UAC99/U206/B (-2358.5 , 285.5)
*       1805 = UAC99/F6 (-2354.5 , 314)
*       1805 = UAC98/F (-2311.5 , 294)
*       1805 = UAC98/U206/B (-1988 , 285.5)
*       1805 = UAC98/F6 (-1984 , 314)
*       1805 = UAC97/F (-1947.5 , 294)
*       1805 = UAC97/U206/B (-1624 , 285.5)
*       1805 = UAC97/F6 (-1620 , 314)
*       1805 = UAC96/F (-1579.5 , 294)
*       1805 = UAC96/U206/B (-1256 , 285.5)
*       1805 = UAC96/F6 (-1252 , 314)
*       1805 = UAC62/F (-1208 , 294)
*       1805 = UAC63/F (-844.5 , 294)
*       1805 = UAC62/U206/B (-884.5 , 285.5)
*       1805 = UAC62/F6 (-880.5 , 314)
*       1805 = UAC63/U206/B (-521 , 285.5)
*       1805 = UAC63/F6 (-517 , 314)
*       1805 = UAC64/F (-480 , 294)
*       1805 = UAC65/F (-116.5 , 294)
*       1805 = UAC64/U206/B (-156.5 , 285.5)
*       1805 = UAC64/F6 (-152.5 , 314)
*       1805 = UAC65/U206/B (207 , 285.5)
*       1805 = UAC65/F6 (211 , 314)
*       1812 = UAC62/U222/B (-1015 , 285.5)
*       1812 = UAC62/U206/A (-958 , 290.5)
*       1812 = UAC62/A6 (-956.5 , 320)
*       1812 = UAC66/S (-848 , 364)
*       1812 = UAC66/U218/Vout (-682.5 , 416)
*       1813 = UAC62/U222/Vout (-1053 , 297.5)
*       1813 = UAC62/U218/A (-1082 , 246.5)
*       1820 = UAC62/U219/OUT (-1156.5 , 274)
*       1820 = UAC62/U262/vin (-1106.5 , 286)
*       1821 = UAC62/U262/vout (-1121 , 287.5)
*       1821 = UAC62/U222/A (-1088.5 , 290.5)
*       1822 = UAC62/U238/B (-1144 , 241.5)
*       1822 = UAC62/U220/A (-998.5 , 285.5)
*       1822 = UAC62/C6 (-998.5 , 317.5)
*       1822 = UAC63/U254/Vout (-676 , 199)
*       1822 = UAC63/P (-675 , 172)
*       1822 = UAC62/U236/B (-873 , 241.5)
*       1822 = UAC62/C (-832.5 , 268.5)
*       1823 = UAC62/U245/Vout (-1103.5 , 243)
*       1823 = UAC62/U253/A (-1009.5 , 187.5)
*       1829 = UAC96/U229/Vin (-1355 , 243)
*       1829 = UAC96/U220/OUT (-1356.5 , 274)
*       1834 = UAC96/U206/Vout (-1294 , 297.5)
*       1834 = UAC96/U236/A (-1271 , 241.5)
*       1834 = UAC96/U235/B (-1289 , 241.5)
*       1843 = UAC96/U222/Vout (-1424.5 , 297.5)
*       1843 = UAC96/U218/A (-1453.5 , 246.5)
*       1845 = UAC96/U218/B (-1380 , 241.5)
*       1845 = UAC96/U229/Vout (-1341 , 243)
*       1851 = UAC96/U206/A (-1329.5 , 290.5)
*       1851 = UAC96/A6 (-1328 , 320)
*       1851 = UAC96/U222/B (-1386.5 , 285.5)
*       1851 = UAC59/S (-1211.5 , 364)
*       1851 = UAC59/U218/Vout (-1046 , 416)
*       1852 = UAC96/U219/OUT (-1528 , 274)
*       1852 = UAC96/U262/vin (-1478 , 286)
*       1853 = UAC96/U262/vout (-1492.5 , 287.5)
*       1853 = UAC96/U222/A (-1460 , 290.5)
*       1854 = UAC96/U238/B (-1515.5 , 241.5)
*       1854 = UAC96/U220/A (-1370 , 285.5)
*       1854 = UAC96/C6 (-1370 , 317.5)
*       1854 = UAC62/U254/Vout (-1039.5 , 199)
*       1854 = UAC62/P (-1038.5 , 172)
*       1854 = UAC96/U236/B (-1244.5 , 241.5)
*       1854 = UAC96/C (-1204 , 268.5)
*       1860 = UAC97/U206/Vout (-1662 , 297.5)
*       1860 = UAC97/U236/A (-1639 , 241.5)
*       1860 = UAC97/U235/B (-1657 , 241.5)
*       1867 = UAC97/U206/A (-1697.5 , 290.5)
*       1867 = UAC97/A6 (-1696 , 320)
*       1867 = UAC97/U222/B (-1754.5 , 285.5)
*       1867 = UAC91/S (-1583 , 364)
*       1867 = UAC91/U218/Vout (-1417.5 , 416)
*       1868 = UAC97/U229/Vin (-1723 , 243)
*       1868 = UAC97/U220/OUT (-1724.5 , 274)
*       1877 = UAC97/U262/vout (-1860.5 , 287.5)
*       1877 = UAC97/U222/A (-1828 , 290.5)
*       1880 = UAC97/U218/A (-1821.5 , 246.5)
*       1880 = UAC97/U222/Vout (-1792.5 , 297.5)
*       1883 = UAC97/U219/OUT (-1896 , 274)
*       1883 = UAC97/U262/vin (-1846 , 286)
*       1886 = UAC97/U238/B (-1883.5 , 241.5)
*       1886 = UAC97/U220/A (-1738 , 285.5)
*       1886 = UAC97/C6 (-1738 , 317.5)
*       1886 = UAC97/U236/B (-1612.5 , 241.5)
*       1886 = UAC96/U254/Vout (-1411 , 199)
*       1886 = UAC96/P (-1410 , 172)
*       1886 = UAC97/C (-1572 , 268.5)
*       1890 = UAC98/U206/Vout (-2026 , 297.5)
*       1890 = UAC98/U236/A (-2003 , 241.5)
*       1890 = UAC98/U235/B (-2021 , 241.5)
*       1892 = UAC98/U238/B (-2247.5 , 241.5)
*       1892 = UAC98/U220/A (-2102 , 285.5)
*       1892 = UAC98/C6 (-2102 , 317.5)
*       1892 = UAC97/U254/Vout (-1779 , 199)
*       1892 = UAC97/P (-1778 , 172)
*       1892 = UAC98/U236/B (-1976.5 , 241.5)
*       1892 = UAC98/C (-1936 , 268.5)
*       1895 = UAC98/U246/Vin (-1995 , 199)
*       1895 = UAC98/U236/OUT (-1989.5 , 230)
*       1904 = UAC98/U222/B (-2118.5 , 285.5)
*       1904 = UAC98/U206/A (-2061.5 , 290.5)
*       1904 = UAC98/A6 (-2060 , 320)
*       1904 = UAC92/S (-1951 , 364)
*       1904 = UAC92/U218/Vout (-1785.5 , 416)
*       1905 = UAC98/U222/Vout (-2156.5 , 297.5)
*       1905 = UAC98/U218/A (-2185.5 , 246.5)
*       1911 = UAC98/U229/Vin (-2087 , 243)
*       1911 = UAC98/U220/OUT (-2088.5 , 274)
*       1914 = UAC98/U219/OUT (-2260 , 274)
*       1914 = UAC98/U262/vin (-2210 , 286)
*       1915 = UAC98/U262/vout (-2224.5 , 287.5)
*       1915 = UAC98/U222/A (-2192 , 290.5)
*       1916 = UAC98/U245/Vout (-2207 , 243)
*       1916 = UAC98/U253/A (-2113 , 187.5)
*       1922 = UAC99/U229/Vin (-2457.5 , 243)
*       1922 = UAC99/U220/OUT (-2459 , 274)
*       1925 = UAC99/U206/Vout (-2396.5 , 297.5)
*       1925 = UAC99/U235/B (-2391.5 , 241.5)
*       1925 = UAC99/U236/A (-2373.5 , 241.5)
*       1933 = UAC99/U206/A (-2432 , 290.5)
*       1933 = UAC99/A6 (-2430.5 , 320)
*       1933 = UAC99/U222/B (-2489 , 285.5)
*       1933 = UAC93/S (-2315 , 364)
*       1933 = UAC93/U218/Vout (-2149.5 , 416)
*       1937 = UAC99/U222/Vout (-2527 , 297.5)
*       1937 = UAC99/U218/A (-2556 , 246.5)
*       1939 = UAC99/U218/B (-2482.5 , 241.5)
*       1939 = UAC99/U229/Vout (-2443.5 , 243)
*       1945 = UAC99/U262/vout (-2595 , 287.5)
*       1945 = UAC99/U222/A (-2562.5 , 290.5)
*       1946 = UAC99/U238/B (-2618 , 241.5)
*       1946 = UAC99/U220/A (-2472.5 , 285.5)
*       1946 = UAC99/C6 (-2472.5 , 317.5)
*       1946 = UAC98/U254/Vout (-2143 , 199)
*       1946 = UAC98/P (-2142 , 172)
*       1946 = UAC99/U236/B (-2347 , 241.5)
*       1946 = UAC99/C (-2306.5 , 268.5)
*       1949 = UAC99/U219/OUT (-2630.5 , 274)
*       1949 = UAC99/U262/vin (-2580.5 , 286)
*       1953 = UAC100/U206/Vout (-2763.5 , 297.5)
*       1953 = UAC100/U236/A (-2740.5 , 241.5)
*       1953 = UAC100/U235/B (-2758.5 , 241.5)
*       1959 = UAC100/U206/A (-2799 , 290.5)
*       1959 = UAC100/A6 (-2797.5 , 320)
*       1959 = UAC100/U222/B (-2856 , 285.5)
*       1959 = UAC94/S (-2685.5 , 364)
*       1959 = UAC94/U218/Vout (-2520 , 416)
*       1960 = UAC100/U229/Vin (-2824.5 , 243)
*       1960 = UAC100/U220/OUT (-2826 , 274)
*       1968 = UAC100/U262/vout (-2962 , 287.5)
*       1968 = UAC100/U222/A (-2929.5 , 290.5)
*       1973 = UAC100/U218/A (-2923 , 246.5)
*       1973 = UAC100/U222/Vout (-2894 , 297.5)
*       1976 = UAC100/U238/B (-2985 , 241.5)
*       1976 = UAC100/U220/A (-2839.5 , 285.5)
*       1976 = UAC100/C6 (-2839.5 , 317.5)
*       1976 = UAC100/U236/B (-2714 , 241.5)
*       1976 = UAC99/U254/Vout (-2513.5 , 199)
*       1976 = UAC99/P (-2512.5 , 172)
*       1976 = UAC100/C (-2673.5 , 268.5)
*       1977 = UAC100/U219/OUT (-2997.5 , 274)
*       1977 = UAC100/U262/vin (-2947.5 , 286)
*       1983 = UAC101/U206/Vout (-3135 , 297.5)
*       1983 = UAC101/U236/A (-3112 , 241.5)
*       1983 = UAC101/U235/B (-3130 , 241.5)
*       1994 = UAC101/U222/B (-3227.5 , 285.5)
*       1994 = UAC101/U206/A (-3170.5 , 290.5)
*       1994 = UAC101/A6 (-3169 , 320)
*       1994 = UAC95/S (-3052.5 , 364)
*       1994 = UAC95/U218/Vout (-2887 , 416)
*       1995 = UAC101/U229/Vin (-3196 , 243)
*       1995 = UAC101/U220/OUT (-3197.5 , 274)
*       2003 = UAC101/U219/OUT (-3369 , 274)
*       2003 = UAC101/U262/vin (-3319 , 286)
*       2004 = UAC101/U262/vout (-3333.5 , 287.5)
*       2004 = UAC101/U222/A (-3301 , 290.5)
*       2005 = UAC101/U238/B (-3356.5 , 241.5)
*       2005 = UAC101/U220/A (-3211 , 285.5)
*       2005 = UAC101/C6 (-3211 , 317.5)
*       2005 = UAC100/U254/Vout (-2880.5 , 199)
*       2005 = UAC100/P (-2879.5 , 172)
*       2005 = UAC101/U236/B (-3085.5 , 241.5)
*       2005 = UAC101/C (-3045 , 268.5)
*       2006 = UAC101/U245/Vout (-3316 , 243)
*       2006 = UAC101/U253/A (-3222 , 187.5)
*       2007 = UAC101/U218/A (-3294.5 , 246.5)
*       2007 = UAC101/U222/Vout (-3265.5 , 297.5)
*       2011 = UAC120/U228/vin (-3635.5 , 285.5)
*       2011 = UAC120/U227/O/P (-3651 , 293.5)
*       2014 = UAC120/U223/vin (-3727.5 , 285.5)
*       2014 = UAC120/U222/OUT (-3758 , 274)
*       2017 = UAC120/Fn (-3810 , 251.5)
*       2017 = UAC120/U229/B (-3632 , 240)
*       2017 = UAC120/F (-3628.5 , 325.5)
*       2017 = Q2 (-3681.5 , 360.5)
*       2017 = UAC119/Qn (-3444.5 , 360.5)
*       2017 = UAC119/U220/Vout (-3279 , 369.5)
*       2018 = UAC65/U253/C (122 , 187.5)
*       2018 = UAC65/U247/Vout (166 , 199)
*       2019 = UAC65/U247/Vin (152 , 199)
*       2019 = UAC65/U235/OUT (161 , 230)
*       2020 = UAC65/U246/Vin (200 , 199)
*       2020 = UAC65/U236/OUT (205.5 , 230)
*       2023 = UAC65/U218/B (83 , 241.5)
*       2023 = UAC65/U229/Vout (122 , 243)
*       2024 = UAC65/U254/Vin (38 , 199)
*       2024 = UAC65/U253/OUT (72.5 , 187.5)
*       2025 = UAC65/U253/B (94.5 , 188)
*       2025 = UAC65/U246/Vout (214 , 199)
*       2030 = UAC70/U262/vout (-30 , 126)
*       2030 = UAC70/U222/A (2.5 , 129)
*       2031 = UAC65/U245/Vin (-26 , 243)
*       2031 = UAC65/U238/OUT (-65.5 , 230)
*       2032 = UAC64/U246/Vin (-163.5 , 199)
*       2032 = UAC64/U236/OUT (-158 , 230)
*       2034 = UAC64/U253/B (-269 , 188)
*       2034 = UAC64/U246/Vout (-149.5 , 199)
*       2035 = UAC64/U253/C (-241.5 , 187.5)
*       2035 = UAC64/U247/Vout (-197.5 , 199)
*       2036 = UAC64/U247/Vin (-211.5 , 199)
*       2036 = UAC64/U235/OUT (-202.5 , 230)
*       2039 = UAC69/U206/Vout (-195 , 136)
*       2039 = UAC69/U236/A (-172 , 80)
*       2039 = UAC69/U235/B (-190 , 80)
*       2041 = UAC64/U253/OUT (-291 , 187.5)
*       2041 = UAC64/U254/Vin (-325.5 , 199)
*       2042 = UAC64/U253/A (-281.5 , 187.5)
*       2042 = UAC64/U245/Vout (-375.5 , 243)
*       2045 = UAC64/U238/OUT (-429 , 230)
*       2045 = UAC64/U245/Vin (-389.5 , 243)
*       2046 = UAC63/U247/Vin (-576 , 199)
*       2046 = UAC63/U235/OUT (-567 , 230)
*       2047 = UAC63/U246/Vin (-528 , 199)
*       2047 = UAC63/U236/OUT (-522.5 , 230)
*       2050 = UAC63/U218/B (-645 , 241.5)
*       2050 = UAC63/U229/Vout (-606 , 243)
*       2051 = UAC63/U253/B (-633.5 , 188)
*       2051 = UAC63/U246/Vout (-514 , 199)
*       2052 = UAC63/U253/C (-606 , 187.5)
*       2052 = UAC63/U247/Vout (-562 , 199)
*       2056 = UAC63/U253/A (-646 , 187.5)
*       2056 = UAC63/U245/Vout (-740 , 243)
*       2057 = UAC63/U254/Vin (-690 , 199)
*       2057 = UAC63/U253/OUT (-655.5 , 187.5)
*       2058 = UAC68/U218/A (-719 , 85)
*       2058 = UAC68/U222/Vout (-690 , 136)
*       2060 = UAC63/U238/OUT (-793.5 , 230)
*       2060 = UAC63/U245/Vin (-754 , 243)
*       2061 = UAC62/U253/C (-969.5 , 187.5)
*       2061 = UAC62/U247/Vout (-925.5 , 199)
*       2062 = UAC62/U247/Vin (-939.5 , 199)
*       2062 = UAC62/U235/OUT (-930.5 , 230)
*       2063 = UAC62/U246/Vin (-891.5 , 199)
*       2063 = UAC62/U236/OUT (-886 , 230)
*       2067 = UAC62/U218/B (-1008.5 , 241.5)
*       2067 = UAC62/U229/Vout (-969.5 , 243)
*       2068 = UAC62/U254/Vin (-1053.5 , 199)
*       2068 = UAC62/U253/OUT (-1019 , 187.5)
*       2069 = UAC62/U253/B (-997 , 188)
*       2069 = UAC62/U246/Vout (-877.5 , 199)
*       2073 = UAC62/U245/Vin (-1117.5 , 243)
*       2073 = UAC62/U238/OUT (-1157 , 230)
*       2074 = UAC121/U220/B (-3917 , 33.5)
*       2074 = UAC121/U230/vout (-3897 , 77.5)
*       2074 = UAC121/Fn (-3881 , 101.5)
*       2074 = UAC109/F (-3787 , 132.5)
*       2074 = UAC109/U206/B (-3463.5 , 124)
*       2074 = UAC109/F6 (-3459.5 , 152.5)
*       2074 = UAC107/F (-3414.5 , 132.5)
*       2074 = UAC107/U206/B (-3091 , 124)
*       2074 = UAC107/F6 (-3087 , 152.5)
*       2074 = UAC106/F (-3043 , 132.5)
*       2074 = UAC106/U206/B (-2719.5 , 124)
*       2074 = UAC106/F6 (-2715.5 , 152.5)
*       2074 = UAC105/F (-2676 , 132.5)
*       2074 = UAC105/U206/B (-2352.5 , 124)
*       2074 = UAC105/F6 (-2348.5 , 152.5)
*       2074 = UAC104/F (-2305.5 , 132.5)
*       2074 = UAC104/U206/B (-1982 , 124)
*       2074 = UAC104/F6 (-1978 , 152.5)
*       2074 = UAC103/F (-1941.5 , 132.5)
*       2074 = UAC103/U206/B (-1618 , 124)
*       2074 = UAC103/F6 (-1614 , 152.5)
*       2074 = UAC102/F (-1573.5 , 132.5)
*       2074 = UAC102/U206/B (-1250 , 124)
*       2074 = UAC67/F (-1208.5 , 132.5)
*       2074 = UAC102/F6 (-1246 , 152.5)
*       2074 = UAC67/U206/B (-885 , 124)
*       2074 = UAC67/F6 (-881 , 152.5)
*       2074 = UAC68/F (-845 , 132.5)
*       2074 = UAC68/U206/B (-521.5 , 124)
*       2074 = UAC68/F6 (-517.5 , 152.5)
*       2074 = UAC69/F (-480.5 , 132.5)
*       2074 = UAC69/U206/B (-157 , 124)
*       2074 = UAC70/F (-117 , 132.5)
*       2074 = UAC69/F6 (-153 , 152.5)
*       2074 = UAC70/U206/B (206.5 , 124)
*       2074 = UAC70/F6 (210.5 , 152.5)
*       2075 = UAC96/U246/Vin (-1263 , 199)
*       2075 = UAC96/U236/OUT (-1257.5 , 230)
*       2077 = UAC96/U253/B (-1368.5 , 188)
*       2077 = UAC96/U246/Vout (-1249 , 199)
*       2078 = UAC96/U253/C (-1341 , 187.5)
*       2078 = UAC96/U247/Vout (-1297 , 199)
*       2079 = UAC96/U247/Vin (-1311 , 199)
*       2079 = UAC96/U235/OUT (-1302 , 230)
*       2084 = UAC96/U253/A (-1381 , 187.5)
*       2084 = UAC96/U245/Vout (-1475 , 243)
*       2085 = UAC96/U254/Vin (-1425 , 199)
*       2085 = UAC96/U253/OUT (-1390.5 , 187.5)
*       2088 = UAC96/U238/OUT (-1528.5 , 230)
*       2088 = UAC96/U245/Vin (-1489 , 243)
*       2089 = UAC97/U247/Vin (-1679 , 199)
*       2089 = UAC97/U235/OUT (-1670 , 230)
*       2090 = UAC97/U246/Vin (-1631 , 199)
*       2090 = UAC97/U236/OUT (-1625.5 , 230)
*       2093 = UAC97/U218/B (-1748 , 241.5)
*       2093 = UAC97/U229/Vout (-1709 , 243)
*       2094 = UAC97/U253/B (-1736.5 , 188)
*       2094 = UAC97/U246/Vout (-1617 , 199)
*       2095 = UAC97/U253/C (-1709 , 187.5)
*       2095 = UAC97/U247/Vout (-1665 , 199)
*       2099 = UAC97/U253/A (-1749 , 187.5)
*       2099 = UAC97/U245/Vout (-1843 , 243)
*       2100 = UAC97/U254/Vin (-1793 , 199)
*       2100 = UAC97/U253/OUT (-1758.5 , 187.5)
*       2102 = UAC97/U238/OUT (-1896.5 , 230)
*       2102 = UAC97/U245/Vin (-1857 , 243)
*       2103 = UAC98/U253/C (-2073 , 187.5)
*       2103 = UAC98/U247/Vout (-2029 , 199)
*       2104 = UAC98/U247/Vin (-2043 , 199)
*       2104 = UAC98/U235/OUT (-2034 , 230)
*       2107 = UAC104/U238/B (-2241.5 , 80)
*       2107 = UAC104/U220/A (-2096 , 124)
*       2107 = UAC104/C6 (-2096 , 156)
*       2107 = UAC103/P (-1772 , 10.5)
*       2107 = UAC104/U236/B (-1970.5 , 80)
*       2107 = UAC104/C (-1930 , 107)
*       2107 = UAC103/U254/Vout (-1773 , 37.5)
*       2108 = UAC98/U218/B (-2112 , 241.5)
*       2108 = UAC98/U229/Vout (-2073 , 243)
*       2109 = UAC98/U254/Vin (-2157 , 199)
*       2109 = UAC98/U253/OUT (-2122.5 , 187.5)
*       2110 = UAC98/U253/B (-2100.5 , 188)
*       2110 = UAC98/U246/Vout (-1981 , 199)
*       2115 = UAC98/U245/Vin (-2221 , 243)
*       2115 = UAC98/U238/OUT (-2260.5 , 230)
*       2116 = UAC99/U246/Vin (-2365.5 , 199)
*       2116 = UAC99/U236/OUT (-2360 , 230)
*       2118 = UAC99/U253/B (-2471 , 188)
*       2118 = UAC99/U246/Vout (-2351.5 , 199)
*       2119 = UAC99/U253/C (-2443.5 , 187.5)
*       2119 = UAC99/U247/Vout (-2399.5 , 199)
*       2120 = UAC99/U247/Vin (-2413.5 , 199)
*       2120 = UAC99/U235/OUT (-2404.5 , 230)
*       2123 = UAC105/U236/A (-2367.5 , 80)
*       2123 = UAC105/U235/B (-2385.5 , 80)
*       2123 = UAC105/U206/Vout (-2390.5 , 136)
*       2125 = UAC99/U253/A (-2483.5 , 187.5)
*       2125 = UAC99/U245/Vout (-2577.5 , 243)
*       2126 = UAC99/U254/Vin (-2527.5 , 199)
*       2126 = UAC99/U253/OUT (-2493 , 187.5)
*       2129 = UAC99/U245/Vin (-2591.5 , 243)
*       2129 = UAC99/U238/OUT (-2631 , 230)
*       2130 = UAC105/U262/vout (-2589 , 126)
*       2130 = UAC105/U222/A (-2556.5 , 129)
*       2131 = UAC100/U247/Vin (-2780.5 , 199)
*       2131 = UAC100/U235/OUT (-2771.5 , 230)
*       2132 = UAC100/U246/Vin (-2732.5 , 199)
*       2132 = UAC100/U236/OUT (-2727 , 230)
*       2135 = UAC100/U218/B (-2849.5 , 241.5)
*       2135 = UAC100/U229/Vout (-2810.5 , 243)
*       2136 = UAC100/U253/B (-2838 , 188)
*       2136 = UAC100/U246/Vout (-2718.5 , 199)
*       2137 = UAC100/U253/C (-2810.5 , 187.5)
*       2137 = UAC100/U247/Vout (-2766.5 , 199)
*       2141 = UAC100/U253/A (-2850.5 , 187.5)
*       2141 = UAC100/U245/Vout (-2944.5 , 243)
*       2142 = UAC100/U254/Vin (-2894.5 , 199)
*       2142 = UAC100/U253/OUT (-2860 , 187.5)
*       2145 = UAC100/U238/OUT (-2998 , 230)
*       2145 = UAC100/U245/Vin (-2958.5 , 243)
*       2146 = UAC101/U253/C (-3182 , 187.5)
*       2146 = UAC101/U247/Vout (-3138 , 199)
*       2147 = UAC101/U247/Vin (-3152 , 199)
*       2147 = UAC101/U235/OUT (-3143 , 230)
*       2148 = UAC101/U246/Vin (-3104 , 199)
*       2148 = UAC101/U236/OUT (-3098.5 , 230)
*       2151 = UAC101/U218/B (-3221 , 241.5)
*       2151 = UAC101/U229/Vout (-3182 , 243)
*       2152 = UAC101/U254/Vin (-3266 , 199)
*       2152 = UAC101/U253/OUT (-3231.5 , 187.5)
*       2153 = UAC101/U253/B (-3209.5 , 188)
*       2153 = UAC101/U246/Vout (-3090 , 199)
*       2158 = UAC101/U245/Vin (-3330 , 243)
*       2158 = UAC101/U238/OUT (-3369.5 , 230)
*       2164 = UAC120/U230/vin (-3614.5 , 240)
*       2164 = UAC120/U229/OUT (-3645 , 228.5)
*       2165 = UAC109/U222/B (-3594 , 124)
*       2165 = UAC109/U206/A (-3537 , 129)
*       2165 = UAC109/A6 (-3535.5 , 158.5)
*       2165 = UAC101/S (-3424.5 , 201.5)
*       2165 = UAC101/U218/Vout (-3259 , 253.5)
*       2166 = UAC120/U227/B (-3664.5 , 300)
*       2166 = UAC120/U226/vout (-3670 , 239)
*       2172 = UAC120/U231/B (-3737 , 195)
*       2172 = UAC120/Pn (-3737.5 , 168.5)
*       2172 = UAC101/U254/Vout (-3252 , 199)
*       2172 = UAC101/P (-3251 , 172)
*       2173 = UAC120/U232/vin (-3719.5 , 195)
*       2173 = UAC120/U231/OUT (-3750 , 183.5)
*       2174 = UAC120/U226/vin (-3698.5 , 240)
*       2174 = UAC120/U225/OUT (-3729 , 228.5)
*       2175 = UAC120/U220/A (-3679.5 , 200)
*       2175 = UAC120/U232/vout (-3691 , 194)
*       2176 = UAC120/U225/A (-3742.5 , 240)
*       2176 = UAC120/U224/vout (-3754 , 239)
*       2177 = UAC120/U225/B (-3716 , 240)
*       2177 = UAC120/U222/B (-3745 , 285.5)
*       2177 = UAC120/L (-3746 , 323)
*       2177 = Lf1 (-3745.5 , 330.5)
*       2180 = Q1 (-3998.5 , 197.5)
*       2180 = UAC121/Fn (-4121 , 90)
*       2180 = UAC121/U229/B (-3943 , 78.5)
*       2180 = UAC121/F (-3939.5 , 164)
*       2180 = UAC120/Qn (-3809.5 , 198)
*       2180 = UAC120/U220/Vout (-3644 , 207)
*       2183 = UAC70/U236/A (191.5 , 80)
*       2183 = UAC70/U235/B (173.5 , 80)
*       2183 = UAC70/U206/Vout (168.5 , 136)
*       2193 = UAC70/U218/B (82.5 , 80)
*       2193 = UAC70/U229/Vout (121.5 , 81.5)
*       2194 = UAC70/U229/Vin (107.5 , 81.5)
*       2194 = UAC70/U220/OUT (106 , 112.5)
*       2195 = UAC70/U218/A (9 , 85)
*       2195 = UAC70/U222/Vout (38 , 136)
*       2197 = UAC121/U228/vout (-3918 , 123)
*       2197 = UAC121/D (-3881.5 , 118.5)
*       2197 = UAC109/D (-3787 , 120.5)
*       2197 = UAC109/U219/B (-3722.5 , 124)
*       2197 = UAC109/U220/B (-3551 , 124)
*       2197 = UAC107/D (-3414.5 , 120.5)
*       2197 = UAC107/U219/B (-3350 , 124)
*       2197 = UAC107/U220/B (-3178.5 , 124)
*       2197 = UAC106/D (-3043 , 120.5)
*       2197 = UAC106/U219/B (-2978.5 , 124)
*       2197 = UAC106/U220/B (-2807 , 124)
*       2197 = UAC105/D (-2676 , 120.5)
*       2197 = UAC105/U219/B (-2611.5 , 124)
*       2197 = UAC105/U220/B (-2440 , 124)
*       2197 = UAC104/D (-2305.5 , 120.5)
*       2197 = UAC104/U219/B (-2241 , 124)
*       2197 = UAC104/U220/B (-2069.5 , 124)
*       2197 = UAC103/D (-1941.5 , 120.5)
*       2197 = UAC103/U219/B (-1877 , 124)
*       2197 = UAC103/U220/B (-1705.5 , 124)
*       2197 = UAC102/D (-1573.5 , 120.5)
*       2197 = UAC102/U219/B (-1509 , 124)
*       2197 = UAC102/U220/B (-1337.5 , 124)
*       2197 = UAC67/D (-1208.5 , 120.5)
*       2197 = UAC67/U219/B (-1144 , 124)
*       2197 = UAC67/U220/B (-972.5 , 124)
*       2197 = UAC68/D (-845 , 120.5)
*       2197 = UAC68/U219/B (-780.5 , 124)
*       2197 = UAC68/U220/B (-609 , 124)
*       2197 = UAC69/D (-480.5 , 120.5)
*       2197 = UAC69/U219/B (-416 , 124)
*       2197 = UAC69/U220/B (-244.5 , 124)
*       2197 = UAC70/D (-117 , 120.5)
*       2197 = UAC70/U219/B (-52.5 , 124)
*       2197 = UAC70/U220/B (119 , 124)
*       2197 = UAC121/Dn (-3919.5 , 165)
*       2197 = UAC109/D6 (-3723 , 151)
*       2197 = UAC107/D6 (-3350.5 , 151)
*       2197 = UAC106/D6 (-2979 , 151)
*       2197 = UAC105/D6 (-2612 , 151)
*       2197 = UAC104/D6 (-2241.5 , 151)
*       2197 = UAC103/D6 (-1877.5 , 151)
*       2197 = UAC102/D6 (-1509.5 , 151)
*       2197 = UAC67/D6 (-1144.5 , 151)
*       2197 = UAC68/D6 (-781 , 151)
*       2197 = UAC69/D6 (-416.5 , 151)
*       2197 = UAC70/D6 (-53 , 151)
*       2201 = UAC70/U222/B (76 , 124)
*       2201 = UAC121/U223/vout (-4010 , 123)
*       2201 = UAC121/An (-4011 , 167)
*       2201 = UAC70/U206/A (133 , 129)
*       2201 = UAC70/A6 (134.5 , 158.5)
*       2206 = UAC70/U245/Vout (-12.5 , 81.5)
*       2206 = UAC70/U253/A (81.5 , 26)
*       2207 = UAC70/U245/Vin (-26.5 , 81.5)
*       2207 = UAC70/U238/OUT (-66 , 68.5)
*       2208 = UAC70/U262/vin (-15.5 , 124.5)
*       2208 = UAC70/U219/OUT (-65.5 , 112.5)
*       2211 = UAC70/S (-121 , 40)
*       2211 = UAC74/U222/B (75.5 , -38.5)
*       2211 = UAC74/U206/A (132.5 , -33.5)
*       2211 = UAC74/A6 (134 , -4)
*       2211 = UAC70/U218/Vout (44.5 , 92)
*       2215 = UAC69/U229/Vin (-256 , 81.5)
*       2215 = UAC69/U220/OUT (-257.5 , 112.5)
*       2218 = UAC69/U222/B (-287.5 , 124)
*       2218 = UAC69/U206/A (-230.5 , 129)
*       2218 = UAC69/A6 (-229 , 158.5)
*       2218 = UAC65/S (-120.5 , 201.5)
*       2218 = UAC65/U218/Vout (45 , 253.5)
*       2223 = UAC69/U254/Vin (-326 , 37.5)
*       2223 = UAC69/U253/OUT (-291.5 , 26)
*       2229 = UAC69/U245/Vout (-376 , 81.5)
*       2229 = UAC69/U253/A (-282 , 26)
*       2230 = UAC69/U218/A (-354.5 , 85)
*       2230 = UAC69/U222/Vout (-325.5 , 136)
*       2232 = UAC69/U218/B (-281 , 80)
*       2232 = UAC69/U229/Vout (-242 , 81.5)
*       2233 = UAC69/U262/vout (-393.5 , 126)
*       2233 = UAC69/U222/A (-361 , 129)
*       2238 = UAC69/S (-484.5 , 40)
*       2238 = UAC73/U206/A (-231 , -33.5)
*       2238 = UAC73/A6 (-229.5 , -4)
*       2238 = UAC73/U222/B (-288 , -38.5)
*       2238 = UAC69/U218/Vout (-319 , 92)
*       2239 = UAC69/U238/OUT (-429.5 , 68.5)
*       2239 = UAC69/U245/Vin (-390 , 81.5)
*       2240 = UAC69/U238/B (-416.5 , 80)
*       2240 = UAC69/U220/A (-271 , 124)
*       2240 = UAC69/C6 (-271 , 156)
*       2240 = UAC70/P (52.5 , 10.5)
*       2240 = UAC69/U236/B (-145.5 , 80)
*       2240 = UAC69/C (-105 , 107)
*       2240 = UAC70/U254/Vout (51.5 , 37.5)
*       2241 = UAC69/U219/OUT (-429 , 112.5)
*       2241 = UAC69/U262/vin (-379 , 124.5)
*       2246 = UAC68/U236/A (-536.5 , 80)
*       2246 = UAC68/U235/B (-554.5 , 80)
*       2246 = UAC68/U206/Vout (-559.5 , 136)
*       2252 = UAC68/U218/B (-645.5 , 80)
*       2252 = UAC68/U229/Vout (-606.5 , 81.5)
*       2253 = UAC68/U229/Vin (-620.5 , 81.5)
*       2253 = UAC68/U220/OUT (-622 , 112.5)
*       2257 = UAC68/U222/B (-652 , 124)
*       2257 = UAC68/U206/A (-595 , 129)
*       2257 = UAC68/A6 (-593.5 , 158.5)
*       2257 = UAC64/S (-484 , 201.5)
*       2257 = UAC64/U218/Vout (-318.5 , 253.5)
*       2266 = UAC68/U245/Vout (-740.5 , 81.5)
*       2266 = UAC68/U253/A (-646.5 , 26)
*       2267 = UAC68/U254/Vin (-690.5 , 37.5)
*       2267 = UAC68/U253/OUT (-656 , 26)
*       2268 = UAC68/U262/vout (-758 , 126)
*       2268 = UAC68/U222/A (-725.5 , 129)
*       2270 = UAC68/S (-849 , 40)
*       2270 = UAC72/U206/A (-595.5 , -33.5)
*       2270 = UAC72/A6 (-594 , -4)
*       2270 = UAC72/U222/B (-652.5 , -38.5)
*       2270 = UAC68/U218/Vout (-683.5 , 92)
*       2271 = UAC68/U238/OUT (-794 , 68.5)
*       2271 = UAC68/U245/Vin (-754.5 , 81.5)
*       2272 = UAC68/U219/OUT (-793.5 , 112.5)
*       2272 = UAC68/U262/vin (-743.5 , 124.5)
*       2274 = UAC68/U238/B (-781 , 80)
*       2274 = UAC68/U220/A (-635.5 , 124)
*       2274 = UAC68/C6 (-635.5 , 156)
*       2274 = UAC68/U236/B (-510 , 80)
*       2274 = UAC69/P (-311 , 10.5)
*       2274 = UAC68/C (-469.5 , 107)
*       2274 = UAC69/U254/Vout (-312 , 37.5)
*       2279 = UAC67/U236/A (-900 , 80)
*       2279 = UAC67/U235/B (-918 , 80)
*       2279 = UAC67/U206/Vout (-923 , 136)
*       2280 = UAC67/U229/Vin (-984 , 81.5)
*       2280 = UAC67/U220/OUT (-985.5 , 112.5)
*       2291 = UAC67/U218/B (-1009 , 80)
*       2291 = UAC67/U229/Vout (-970 , 81.5)
*       2292 = UAC67/U218/A (-1082.5 , 85)
*       2292 = UAC67/U222/Vout (-1053.5 , 136)
*       2294 = UAC67/U262/vout (-1121.5 , 126)
*       2294 = UAC67/U222/A (-1089 , 129)
*       2297 = UAC67/U222/B (-1015.5 , 124)
*       2297 = UAC67/U206/A (-958.5 , 129)
*       2297 = UAC67/A6 (-957 , 158.5)
*       2297 = UAC63/S (-848.5 , 201.5)
*       2297 = UAC63/U218/Vout (-683 , 253.5)
*       2300 = UAC67/U253/B (-997.5 , 26.5)
*       2300 = UAC67/U246/Vout (-878 , 37.5)
*       2302 = UAC67/U245/Vout (-1104 , 81.5)
*       2302 = UAC67/U253/A (-1010 , 26)
*       2303 = UAC67/U245/Vin (-1118 , 81.5)
*       2303 = UAC67/U238/OUT (-1157.5 , 68.5)
*       2304 = UAC67/U262/vin (-1107 , 124.5)
*       2304 = UAC67/U219/OUT (-1157 , 112.5)
*       2305 = UAC67/U238/B (-1144.5 , 80)
*       2305 = UAC67/U220/A (-999 , 124)
*       2305 = UAC67/C6 (-999 , 156)
*       2305 = UAC68/P (-675.5 , 10.5)
*       2305 = UAC67/U236/B (-873.5 , 80)
*       2305 = UAC67/C (-833 , 107)
*       2305 = UAC68/U254/Vout (-676.5 , 37.5)
*       2308 = UAC67/S (-1212.5 , 40)
*       2308 = UAC71/U222/B (-1016 , -38.5)
*       2308 = UAC71/U206/A (-959 , -33.5)
*       2308 = UAC71/A6 (-957.5 , -4)
*       2308 = UAC67/U218/Vout (-1047 , 92)
*       2313 = UAC102/U253/C (-1335 , 26)
*       2313 = UAC102/U247/Vout (-1291 , 37.5)
*       2314 = UAC102/U229/Vin (-1349 , 81.5)
*       2314 = UAC102/U220/OUT (-1350.5 , 112.5)
*       2317 = UAC102/U236/A (-1265 , 80)
*       2317 = UAC102/U235/B (-1283 , 80)
*       2317 = UAC102/U206/Vout (-1288 , 136)
*       2324 = UAC102/U245/Vout (-1469 , 81.5)
*       2324 = UAC102/U253/A (-1375 , 26)
*       2325 = UAC102/U218/A (-1447.5 , 85)
*       2325 = UAC102/U222/Vout (-1418.5 , 136)
*       2327 = UAC102/U218/B (-1374 , 80)
*       2327 = UAC102/U229/Vout (-1335 , 81.5)
*       2328 = UAC102/U262/vout (-1486.5 , 126)
*       2328 = UAC102/U222/A (-1454 , 129)
*       2331 = UAC102/U222/B (-1380.5 , 124)
*       2331 = UAC102/U206/A (-1323.5 , 129)
*       2331 = UAC102/A6 (-1322 , 158.5)
*       2331 = UAC62/S (-1212 , 201.5)
*       2331 = UAC62/U218/Vout (-1046.5 , 253.5)
*       2335 = UAC102/S (-1577.5 , 40)
*       2335 = Sf4 (-1575.5 , 40.5)
*       2335 = UAC102/U218/Vout (-1412 , 92)
*       2336 = UAC102/U238/OUT (-1522.5 , 68.5)
*       2336 = UAC102/U245/Vin (-1483 , 81.5)
*       2337 = UAC102/U238/B (-1509.5 , 80)
*       2337 = UAC102/U220/A (-1364 , 124)
*       2337 = UAC102/C6 (-1364 , 156)
*       2337 = UAC67/P (-1039 , 10.5)
*       2337 = UAC102/U236/B (-1238.5 , 80)
*       2337 = UAC102/C (-1198 , 107)
*       2337 = UAC67/U254/Vout (-1040 , 37.5)
*       2338 = UAC102/U219/OUT (-1522 , 112.5)
*       2338 = UAC102/U262/vin (-1472 , 124.5)
*       2343 = UAC103/U236/A (-1633 , 80)
*       2343 = UAC103/U235/B (-1651 , 80)
*       2343 = UAC103/U206/Vout (-1656 , 136)
*       2350 = UAC103/U218/B (-1742 , 80)
*       2350 = UAC103/U229/Vout (-1703 , 81.5)
*       2351 = UAC103/U229/Vin (-1717 , 81.5)
*       2351 = UAC103/U220/OUT (-1718.5 , 112.5)
*       2355 = UAC103/U222/B (-1748.5 , 124)
*       2355 = UAC103/U206/A (-1691.5 , 129)
*       2355 = UAC103/A6 (-1690 , 158.5)
*       2355 = UAC96/S (-1583.5 , 201.5)
*       2355 = UAC96/U218/Vout (-1418 , 253.5)
*       2364 = UAC103/U245/Vout (-1837 , 81.5)
*       2364 = UAC103/U253/A (-1743 , 26)
*       2365 = UAC103/U262/vin (-1840 , 124.5)
*       2365 = UAC103/U219/OUT (-1890 , 112.5)
*       2366 = UAC103/U218/A (-1815.5 , 85)
*       2366 = UAC103/U222/Vout (-1786.5 , 136)
*       2367 = UAC103/U262/vout (-1854.5 , 126)
*       2367 = UAC103/U222/A (-1822 , 129)
*       2368 = UAC103/S (-1945.5 , 40)
*       2368 = Sf5 (-1943.5 , 40.5)
*       2368 = UAC103/U218/Vout (-1780 , 92)
*       2369 = UAC103/U245/Vin (-1851 , 81.5)
*       2369 = UAC103/U238/OUT (-1890.5 , 68.5)
*       2371 = UAC103/U238/B (-1877.5 , 80)
*       2371 = UAC103/U220/A (-1732 , 124)
*       2371 = UAC103/C6 (-1732 , 156)
*       2371 = UAC103/U236/B (-1606.5 , 80)
*       2371 = UAC102/P (-1404 , 10.5)
*       2371 = UAC103/C (-1566 , 107)
*       2371 = UAC102/U254/Vout (-1405 , 37.5)
*       2376 = UAC104/U236/A (-1997 , 80)
*       2376 = UAC104/U235/B (-2015 , 80)
*       2376 = UAC104/U206/Vout (-2020 , 136)
*       2377 = UAC104/U229/Vin (-2081 , 81.5)
*       2377 = UAC104/U220/OUT (-2082.5 , 112.5)
*       2388 = UAC104/U218/B (-2106 , 80)
*       2388 = UAC104/U229/Vout (-2067 , 81.5)
*       2389 = UAC104/U218/A (-2179.5 , 85)
*       2389 = UAC104/U222/Vout (-2150.5 , 136)
*       2391 = UAC104/U262/vout (-2218.5 , 126)
*       2391 = UAC104/U222/A (-2186 , 129)
*       2394 = UAC104/U222/B (-2112.5 , 124)
*       2394 = UAC104/U206/A (-2055.5 , 129)
*       2394 = UAC104/A6 (-2054 , 158.5)
*       2394 = UAC97/S (-1951.5 , 201.5)
*       2394 = UAC97/U218/Vout (-1786 , 253.5)
*       2398 = UAC104/U245/Vout (-2201 , 81.5)
*       2398 = UAC104/U253/A (-2107 , 26)
*       2399 = UAC104/U245/Vin (-2215 , 81.5)
*       2399 = UAC104/U238/OUT (-2254.5 , 68.5)
*       2400 = UAC104/U262/vin (-2204 , 124.5)
*       2400 = UAC104/U219/OUT (-2254 , 112.5)
*       2403 = UAC104/S (-2309.5 , 40)
*       2403 = Sf6 (-2308 , 40.5)
*       2403 = UAC104/U218/Vout (-2144 , 92)
*       2408 = UAC105/U229/Vin (-2451.5 , 81.5)
*       2408 = UAC105/U220/OUT (-2453 , 112.5)
*       2418 = UAC105/U245/Vout (-2571.5 , 81.5)
*       2418 = UAC105/U253/A (-2477.5 , 26)
*       2419 = UAC105/U218/A (-2550 , 85)
*       2419 = UAC105/U222/Vout (-2521 , 136)
*       2421 = UAC105/U218/B (-2476.5 , 80)
*       2421 = UAC105/U229/Vout (-2437.5 , 81.5)
*       2424 = UAC105/U222/B (-2483 , 124)
*       2424 = UAC105/U206/A (-2426 , 129)
*       2424 = UAC105/A6 (-2424.5 , 158.5)
*       2424 = UAC98/S (-2315.5 , 201.5)
*       2424 = UAC98/U218/Vout (-2150 , 253.5)
*       2428 = UAC105/S (-2680 , 40)
*       2428 = Sf7 (-2678.5 , 40.5)
*       2428 = UAC105/U218/Vout (-2514.5 , 92)
*       2429 = UAC105/U238/OUT (-2625 , 68.5)
*       2429 = UAC105/U245/Vin (-2585.5 , 81.5)
*       2430 = UAC105/U238/B (-2612 , 80)
*       2430 = UAC105/U220/A (-2466.5 , 124)
*       2430 = UAC105/C6 (-2466.5 , 156)
*       2430 = UAC104/P (-2136 , 10.5)
*       2430 = UAC105/U236/B (-2341 , 80)
*       2430 = UAC105/C (-2300.5 , 107)
*       2430 = UAC104/U254/Vout (-2137 , 37.5)
*       2431 = UAC105/U219/OUT (-2624.5 , 112.5)
*       2431 = UAC105/U262/vin (-2574.5 , 124.5)
*       2436 = UAC106/U236/A (-2734.5 , 80)
*       2436 = UAC106/U235/B (-2752.5 , 80)
*       2436 = UAC106/U206/Vout (-2757.5 , 136)
*       2439 = UAC106/U222/B (-2850 , 124)
*       2439 = UAC106/U206/A (-2793 , 129)
*       2439 = UAC106/A6 (-2791.5 , 158.5)
*       2439 = UAC99/S (-2686 , 201.5)
*       2439 = UAC99/U218/Vout (-2520.5 , 253.5)
*       2443 = UAC106/U218/B (-2843.5 , 80)
*       2443 = UAC106/U229/Vout (-2804.5 , 81.5)
*       2444 = UAC106/U229/Vin (-2818.5 , 81.5)
*       2444 = UAC106/U220/OUT (-2820 , 112.5)
*       2456 = UAC106/U245/Vout (-2938.5 , 81.5)
*       2456 = UAC106/U253/A (-2844.5 , 26)
*       2457 = UAC106/U262/vin (-2941.5 , 124.5)
*       2457 = UAC106/U219/OUT (-2991.5 , 112.5)
*       2458 = UAC106/U218/A (-2917 , 85)
*       2458 = UAC106/U222/Vout (-2888 , 136)
*       2459 = UAC106/U262/vout (-2956 , 126)
*       2459 = UAC106/U222/A (-2923.5 , 129)
*       2460 = UAC106/S (-3047 , 40)
*       2460 = Sf8 (-3047.5 , 41)
*       2460 = UAC106/U218/Vout (-2881.5 , 92)
*       2461 = UAC106/U238/OUT (-2992 , 68.5)
*       2461 = UAC106/U245/Vin (-2952.5 , 81.5)
*       2463 = UAC106/U238/B (-2979 , 80)
*       2463 = UAC106/U220/A (-2833.5 , 124)
*       2463 = UAC106/C6 (-2833.5 , 156)
*       2463 = UAC106/U236/B (-2708 , 80)
*       2463 = UAC105/P (-2506.5 , 10.5)
*       2463 = UAC106/C (-2667.5 , 107)
*       2463 = UAC105/U254/Vout (-2507.5 , 37.5)
*       2467 = UAC107/U236/A (-3106 , 80)
*       2467 = UAC107/U235/B (-3124 , 80)
*       2467 = UAC107/U206/Vout (-3129 , 136)
*       2470 = UAC107/U246/Vin (-3098 , 37.5)
*       2470 = UAC107/U236/OUT (-3092.5 , 68.5)
*       2478 = UAC107/U218/B (-3215 , 80)
*       2478 = UAC107/U229/Vout (-3176 , 81.5)
*       2479 = UAC107/U218/A (-3288.5 , 85)
*       2479 = UAC107/U222/Vout (-3259.5 , 136)
*       2480 = UAC107/U220/OUT (-3191.5 , 112.5)
*       2480 = UAC107/U229/Vin (-3190 , 81.5)
*       2485 = UAC107/U222/B (-3221.5 , 124)
*       2485 = UAC107/U206/A (-3164.5 , 129)
*       2485 = UAC107/A6 (-3163 , 158.5)
*       2485 = UAC100/S (-3053 , 201.5)
*       2485 = UAC100/U218/Vout (-2887.5 , 253.5)
*       2486 = UAC107/U254/Vin (-3260 , 37.5)
*       2486 = UAC107/U253/OUT (-3225.5 , 26)
*       2491 = UAC107/U262/vout (-3327.5 , 126)
*       2491 = UAC107/U222/A (-3295 , 129)
*       2492 = UAC107/U245/Vout (-3310 , 81.5)
*       2492 = UAC107/U253/A (-3216 , 26)
*       2493 = UAC107/U245/Vin (-3324 , 81.5)
*       2493 = UAC107/U238/OUT (-3363.5 , 68.5)
*       2494 = UAC107/U262/vin (-3313 , 124.5)
*       2494 = UAC107/U219/OUT (-3363 , 112.5)
*       2495 = UAC107/U238/B (-3350.5 , 80)
*       2495 = UAC107/U220/A (-3205 , 124)
*       2495 = UAC107/C6 (-3205 , 156)
*       2495 = UAC106/P (-2873.5 , 10.5)
*       2495 = UAC107/U236/B (-3079.5 , 80)
*       2495 = UAC107/C (-3039 , 107)
*       2495 = UAC106/U254/Vout (-2874.5 , 37.5)
*       2498 = UAC107/S (-3418.5 , 40)
*       2498 = Sf9 (-3419 , 41.5)
*       2498 = UAC107/U218/Vout (-3253 , 92)
*       2502 = UAC109/U229/Vin (-3562.5 , 81.5)
*       2502 = UAC109/U220/OUT (-3564 , 112.5)
*       2506 = UAC109/U235/B (-3496.5 , 80)
*       2506 = UAC109/U236/A (-3478.5 , 80)
*       2506 = UAC109/U206/Vout (-3501.5 , 136)
*       2515 = UAC109/U218/B (-3587.5 , 80)
*       2515 = UAC109/U229/Vout (-3548.5 , 81.5)
*       2516 = UAC109/U245/Vout (-3682.5 , 81.5)
*       2516 = UAC109/U253/A (-3588.5 , 26)
*       2517 = UAC109/U218/A (-3661 , 85)
*       2517 = UAC109/U222/Vout (-3632 , 136)
*       2519 = UAC109/U262/vout (-3700 , 126)
*       2519 = UAC109/U222/A (-3667.5 , 129)
*       2524 = UAC109/U245/Vin (-3696.5 , 81.5)
*       2524 = UAC109/U238/OUT (-3736 , 68.5)
*       2525 = UAC109/U238/B (-3723 , 80)
*       2525 = UAC109/U220/A (-3577.5 , 124)
*       2525 = UAC109/C6 (-3577.5 , 156)
*       2525 = UAC107/P (-3245 , 10.5)
*       2525 = UAC109/U236/B (-3452 , 80)
*       2525 = UAC109/C (-3411.5 , 107)
*       2525 = UAC107/U254/Vout (-3246 , 37.5)
*       2526 = UAC109/U219/OUT (-3735.5 , 112.5)
*       2526 = UAC109/U262/vin (-3685.5 , 124.5)
*       2529 = UAC109/S (-3791 , 40)
*       2529 = Sf10 (-3790.5 , 41)
*       2529 = UAC109/U218/Vout (-3625.5 , 92)
*       2531 = UAC121/U230/vin (-3925.5 , 78.5)
*       2531 = UAC121/U229/OUT (-3956 , 67)
*       2532 = UAC121/U226/vout (-3981 , 77.5)
*       2532 = UAC121/U227/B (-3975.5 , 138.5)
*       2533 = UAC121/U228/vin (-3946.5 , 124)
*       2533 = UAC121/U227/O/P (-3962 , 132)
*       2538 = UAC121/U226/vin (-4009.5 , 78.5)
*       2538 = UAC121/U225/OUT (-4040 , 67)
*       2539 = UAC121/U225/A (-4053.5 , 78.5)
*       2539 = UAC121/U224/vout (-4065 , 77.5)
*       2540 = UAC121/U225/B (-4027 , 78.5)
*       2540 = UAC121/U222/B (-4056 , 124)
*       2540 = UAC121/L (-4057 , 161.5)
*       2540 = Lf0 (-4056.5 , 165.5)
*       2542 = UAC121/U223/vin (-4038.5 , 124)
*       2542 = UAC121/U222/OUT (-4069 , 112.5)
*       2545 = UAC121/Qn (-4120.5 , 36.5)
*       2545 = UAC126/Vin (-1348 , -37)
*       2545 = UAC121/U220/Vout (-3955 , 45.5)
*       2545 = Q0 (-3952.5 , 56.5)
*       2549 = UAC70/U253/C (121.5 , 26)
*       2549 = UAC70/U247/Vout (165.5 , 37.5)
*       2550 = UAC70/U247/Vin (151.5 , 37.5)
*       2550 = UAC70/U235/OUT (160.5 , 68.5)
*       2551 = UAC70/U246/Vin (199.5 , 37.5)
*       2551 = UAC70/U236/OUT (205 , 68.5)
*       2558 = UAC70/U254/Vin (37.5 , 37.5)
*       2558 = UAC70/U253/OUT (72 , 26)
*       2559 = UAC70/U253/B (94 , 26.5)
*       2559 = UAC70/U246/Vout (213.5 , 37.5)
*       2564 = UAC124/Vout (-1240 , -37)
*       2564 = UAC71/D (-1209 , -42)
*       2564 = UAC71/U219/B (-1144.5 , -38.5)
*       2564 = UAC71/D6 (-1145 , -11.5)
*       2564 = UAC71/U220/B (-973 , -38.5)
*       2564 = UAC72/D (-845.5 , -42)
*       2564 = UAC72/U219/B (-781 , -38.5)
*       2564 = UAC72/D6 (-781.5 , -11.5)
*       2564 = UAC72/U220/B (-609.5 , -38.5)
*       2564 = UAC73/D (-481 , -42)
*       2564 = UAC73/U219/B (-416.5 , -38.5)
*       2564 = UAC73/D6 (-417 , -11.5)
*       2564 = UAC73/U220/B (-245 , -38.5)
*       2564 = UAC74/D (-117.5 , -42)
*       2564 = UAC74/U219/B (-53 , -38.5)
*       2564 = UAC74/D6 (-53.5 , -11.5)
*       2564 = UAC74/U220/B (118.5 , -38.5)
*       2567 = UAC74/U219/OUT (-66 , -50)
*       2567 = UAC74/U262/vin (-16 , -38)
*       2568 = UAC74/U262/vout (-30.5 , -36.5)
*       2568 = UAC74/U222/A (2 , -33.5)
*       2570 = UAC69/U246/Vin (-164 , 37.5)
*       2570 = UAC69/U236/OUT (-158.5 , 68.5)
*       2573 = UAC69/U253/B (-269.5 , 26.5)
*       2573 = UAC69/U246/Vout (-150 , 37.5)
*       2574 = UAC69/U253/C (-242 , 26)
*       2574 = UAC69/U247/Vout (-198 , 37.5)
*       2575 = UAC69/U247/Vin (-212 , 37.5)
*       2575 = UAC69/U235/OUT (-203 , 68.5)
*       2579 = UAC73/U206/Vout (-195.5 , -26.5)
*       2579 = UAC73/U236/A (-172.5 , -82.5)
*       2579 = UAC73/U235/B (-190.5 , -82.5)
*       2587 = UAC73/U218/B (-281.5 , -82.5)
*       2587 = UAC73/U229/Vout (-242.5 , -81)
*       2591 = UAC73/U219/OUT (-429.5 , -50)
*       2591 = UAC73/U262/vin (-379.5 , -38)
*       2592 = UAC73/U262/vout (-394 , -36.5)
*       2592 = UAC73/U222/A (-361.5 , -33.5)
*       2597 = UAC68/U247/Vin (-576.5 , 37.5)
*       2597 = UAC68/U235/OUT (-567.5 , 68.5)
*       2598 = UAC68/U246/Vin (-528.5 , 37.5)
*       2598 = UAC68/U236/OUT (-523 , 68.5)
*       2602 = UAC68/U253/B (-634 , 26.5)
*       2602 = UAC68/U246/Vout (-514.5 , 37.5)
*       2603 = UAC68/U253/C (-606.5 , 26)
*       2603 = UAC68/U247/Vout (-562.5 , 37.5)
*       2611 = UAC72/U262/vout (-758.5 , -36.5)
*       2611 = UAC72/U222/A (-726 , -33.5)
*       2612 = UAC72/U218/A (-719.5 , -77.5)
*       2612 = UAC72/U222/Vout (-690.5 , -26.5)
*       2615 = UAC72/U219/OUT (-794 , -50)
*       2615 = UAC72/U262/vin (-744 , -38)
*       2620 = UAC67/U253/C (-970 , 26)
*       2620 = UAC67/U247/Vout (-926 , 37.5)
*       2621 = UAC67/U247/Vin (-940 , 37.5)
*       2621 = UAC67/U235/OUT (-931 , 68.5)
*       2622 = UAC67/U246/Vin (-892 , 37.5)
*       2622 = UAC67/U236/OUT (-886.5 , 68.5)
*       2630 = UAC67/U254/Vin (-1054 , 37.5)
*       2630 = UAC67/U253/OUT (-1019.5 , 26)
*       2636 = UAC71/U219/OUT (-1157.5 , -50)
*       2636 = UAC71/U262/vin (-1107.5 , -38)
*       2637 = UAC71/U262/vout (-1122 , -36.5)
*       2637 = UAC71/U222/A (-1089.5 , -33.5)
*       2639 = UAC102/U246/Vin (-1257 , 37.5)
*       2639 = UAC102/U236/OUT (-1251.5 , 68.5)
*       2640 = UAC102/U253/B (-1362.5 , 26.5)
*       2640 = UAC102/U246/Vout (-1243 , 37.5)
*       2641 = UAC125/OUT (-1293.5 , -50)
*       2641 = UAC124/Vin (-1254 , -37)
*       2642 = UAC126/Vout (-1334 , -37)
*       2642 = UAC125/A (-1307 , -38.5)
*       2643 = UAC102/U247/Vin (-1305 , 37.5)
*       2643 = UAC102/U235/OUT (-1296 , 68.5)
*       2645 = UAC102/U254/Vin (-1419 , 37.5)
*       2645 = UAC102/U253/OUT (-1384.5 , 26)
*       2646 = UAC103/U247/Vin (-1673 , 37.5)
*       2646 = UAC103/U235/OUT (-1664 , 68.5)
*       2647 = UAC103/U246/Vin (-1625 , 37.5)
*       2647 = UAC103/U236/OUT (-1619.5 , 68.5)
*       2648 = UAC103/U254/Vin (-1787 , 37.5)
*       2648 = UAC103/U253/OUT (-1752.5 , 26)
*       2649 = UAC103/U253/B (-1730.5 , 26.5)
*       2649 = UAC103/U246/Vout (-1611 , 37.5)
*       2650 = UAC103/U253/C (-1703 , 26)
*       2650 = UAC103/U247/Vout (-1659 , 37.5)
*       2651 = UAC104/U246/Vin (-1989 , 37.5)
*       2651 = UAC104/U236/OUT (-1983.5 , 68.5)
*       2652 = UAC104/U253/C (-2067 , 26)
*       2652 = UAC104/U247/Vout (-2023 , 37.5)
*       2653 = UAC104/U247/Vin (-2037 , 37.5)
*       2653 = UAC104/U235/OUT (-2028 , 68.5)
*       2654 = UAC104/U254/Vin (-2151 , 37.5)
*       2654 = UAC104/U253/OUT (-2116.5 , 26)
*       2655 = UAC104/U253/B (-2094.5 , 26.5)
*       2655 = UAC104/U246/Vout (-1975 , 37.5)
*       2656 = UAC105/U246/Vin (-2359.5 , 37.5)
*       2656 = UAC105/U236/OUT (-2354 , 68.5)
*       2657 = UAC105/U253/B (-2465 , 26.5)
*       2657 = UAC105/U246/Vout (-2345.5 , 37.5)
*       2658 = UAC105/U253/C (-2437.5 , 26)
*       2658 = UAC105/U247/Vout (-2393.5 , 37.5)
*       2659 = UAC105/U247/Vin (-2407.5 , 37.5)
*       2659 = UAC105/U235/OUT (-2398.5 , 68.5)
*       2660 = UAC105/U254/Vin (-2521.5 , 37.5)
*       2660 = UAC105/U253/OUT (-2487 , 26)
*       2661 = UAC106/U247/Vin (-2774.5 , 37.5)
*       2661 = UAC106/U235/OUT (-2765.5 , 68.5)
*       2662 = UAC106/U246/Vin (-2726.5 , 37.5)
*       2662 = UAC106/U236/OUT (-2721 , 68.5)
*       2663 = UAC106/U254/Vin (-2888.5 , 37.5)
*       2663 = UAC106/U253/OUT (-2854 , 26)
*       2664 = UAC106/U253/B (-2832 , 26.5)
*       2664 = UAC106/U246/Vout (-2712.5 , 37.5)
*       2665 = UAC106/U253/C (-2804.5 , 26)
*       2665 = UAC106/U247/Vout (-2760.5 , 37.5)
*       2666 = UAC107/U253/C (-3176 , 26)
*       2666 = UAC107/U247/Vout (-3132 , 37.5)
*       2667 = UAC107/U247/Vin (-3146 , 37.5)
*       2667 = UAC107/U235/OUT (-3137 , 68.5)
*       2668 = UAC107/U253/B (-3203.5 , 26.5)
*       2668 = UAC107/U246/Vout (-3084 , 37.5)
*       2669 = UAC109/U246/Vin (-3470.5 , 37.5)
*       2669 = UAC109/U236/OUT (-3465 , 68.5)
*       2670 = UAC109/U253/B (-3576 , 26.5)
*       2670 = UAC109/U246/Vout (-3456.5 , 37.5)
*       2671 = UAC109/U253/C (-3548.5 , 26)
*       2671 = UAC109/U247/Vout (-3504.5 , 37.5)
*       2672 = UAC109/U247/Vin (-3518.5 , 37.5)
*       2672 = UAC109/U235/OUT (-3509.5 , 68.5)
*       2673 = UAC109/U254/Vin (-3632.5 , 37.5)
*       2673 = UAC109/U253/OUT (-3598 , 26)
*       2676 = UAC121/U232/vin (-4030.5 , 33.5)
*       2676 = UAC121/U231/OUT (-4061 , 22)
*       2677 = UAC121/U231/B (-4048 , 33.5)
*       2677 = UAC121/Pn (-4048.5 , 7)
*       2677 = Pf0 (-3887 , 10)
*       2677 = UAC109/P (-3617.5 , 10.5)
*       2677 = UAC109/U254/Vout (-3618.5 , 37.5)
*       2678 = UAC121/U232/vout (-4002 , 32.5)
*       2678 = UAC121/U220/A (-3990.5 , 38.5)
*       2679 = UAC74/U253/C (121 , -136.5)
*       2679 = UAC74/U247/Vout (165 , -125)
*       2680 = UAC74/U247/Vin (151 , -125)
*       2680 = UAC74/U235/OUT (160 , -94)
*       2681 = UAC74/U246/Vin (199 , -125)
*       2681 = UAC74/U236/OUT (204.5 , -94)
*       2682 = UAC74/U236/A (191 , -82.5)
*       2682 = UAC74/U235/B (173 , -82.5)
*       2682 = UAC74/U206/Vout (168 , -26.5)
*       2688 = UAC74/U218/B (82 , -82.5)
*       2688 = UAC74/U229/Vout (121 , -81)
*       2689 = UAC74/U254/Vin (37 , -125)
*       2689 = UAC74/U253/OUT (71.5 , -136.5)
*       2690 = UAC74/U253/B (93.5 , -136)
*       2690 = UAC74/U246/Vout (213 , -125)
*       2691 = UAC74/U229/Vin (107 , -81)
*       2691 = UAC74/U220/OUT (105.5 , -50)
*       2695 = UAC74/U245/Vout (-13 , -81)
*       2695 = UAC74/U253/A (81 , -136.5)
*       2696 = UAC74/U245/Vin (-27 , -81)
*       2696 = UAC74/U238/OUT (-66.5 , -94)
*       2697 = UAC74/U218/A (8.5 , -77.5)
*       2697 = UAC74/U222/Vout (37.5 , -26.5)
*       2699 = UAC74/S (-121.5 , -122.5)
*       2699 = r0 (-131 , -160.5)
*       2699 = UAC74/U218/Vout (44 , -70.5)
*       2700 = UAC73/U246/Vin (-164.5 , -125)
*       2700 = UAC73/U236/OUT (-159 , -94)
*       2702 = UAC73/U253/B (-270 , -136)
*       2702 = UAC73/U246/Vout (-150.5 , -125)
*       2703 = UAC73/U253/C (-242.5 , -136.5)
*       2703 = UAC73/U247/Vout (-198.5 , -125)
*       2704 = UAC73/U247/Vin (-212.5 , -125)
*       2704 = UAC73/U235/OUT (-203.5 , -94)
*       2705 = UAC73/U229/Vin (-256.5 , -81)
*       2705 = UAC73/U220/OUT (-258 , -50)
*       2709 = UAC73/U254/Vin (-326.5 , -125)
*       2709 = UAC73/U253/OUT (-292 , -136.5)
*       2713 = UAC73/U245/Vout (-376.5 , -81)
*       2713 = UAC73/U253/A (-282.5 , -136.5)
*       2714 = UAC73/U218/A (-355 , -77.5)
*       2714 = UAC73/U222/Vout (-326 , -26.5)
*       2716 = UAC73/U238/OUT (-430 , -94)
*       2716 = UAC73/U245/Vin (-390.5 , -81)
*       2717 = UAC73/U238/B (-417 , -82.5)
*       2717 = UAC73/U220/A (-271.5 , -38.5)
*       2717 = UAC73/C6 (-271.5 , -6.5)
*       2717 = UAC74/U254/Vout (51 , -125)
*       2717 = UAC74/P (52 , -152)
*       2717 = UAC73/U236/B (-146 , -82.5)
*       2717 = UAC73/C (-105.5 , -55.5)
*       2719 = UAC72/U247/Vin (-577 , -125)
*       2719 = UAC72/U235/OUT (-568 , -94)
*       2720 = UAC72/U246/Vin (-529 , -125)
*       2720 = UAC72/U236/OUT (-523.5 , -94)
*       2721 = UAC72/U236/A (-537 , -82.5)
*       2721 = UAC72/U235/B (-555 , -82.5)
*       2721 = UAC72/U206/Vout (-560 , -26.5)
*       2722 = r1 (-493.5 , -148)
*       2722 = UAC73/S (-485 , -122.5)
*       2722 = UAC73/U218/Vout (-319.5 , -70.5)
*       2726 = UAC72/U218/B (-646 , -82.5)
*       2726 = UAC72/U229/Vout (-607 , -81)
*       2727 = UAC72/U253/B (-634.5 , -136)
*       2727 = UAC72/U246/Vout (-515 , -125)
*       2728 = UAC72/U253/C (-607 , -136.5)
*       2728 = UAC72/U247/Vout (-563 , -125)
*       2729 = UAC72/U229/Vin (-621 , -81)
*       2729 = UAC72/U220/OUT (-622.5 , -50)
*       2735 = UAC72/U245/Vout (-741 , -81)
*       2735 = UAC72/U253/A (-647 , -136.5)
*       2736 = UAC72/U254/Vin (-691 , -125)
*       2736 = UAC72/U253/OUT (-656.5 , -136.5)
*       2737 = UAC72/S (-849.5 , -122.5)
*       2737 = r2 (-859 , -155)
*       2737 = UAC72/U218/Vout (-684 , -70.5)
*       2738 = UAC72/U238/OUT (-794.5 , -94)
*       2738 = UAC72/U245/Vin (-755 , -81)
*       2740 = UAC72/U238/B (-781.5 , -82.5)
*       2740 = UAC72/U220/A (-636 , -38.5)
*       2740 = UAC72/C6 (-636 , -6.5)
*       2740 = UAC72/U236/B (-510.5 , -82.5)
*       2740 = UAC73/U254/Vout (-312.5 , -125)
*       2740 = UAC73/P (-311.5 , -152)
*       2740 = UAC72/C (-470 , -55.5)
*       2742 = UAC71/U253/C (-970.5 , -136.5)
*       2742 = UAC71/U247/Vout (-926.5 , -125)
*       2743 = UAC71/U247/Vin (-940.5 , -125)
*       2743 = UAC71/U235/OUT (-931.5 , -94)
*       2744 = UAC71/U246/Vin (-892.5 , -125)
*       2744 = UAC71/U236/OUT (-887 , -94)
*       2745 = UAC71/U236/A (-900.5 , -82.5)
*       2745 = UAC71/U235/B (-918.5 , -82.5)
*       2745 = UAC71/U206/Vout (-923.5 , -26.5)
*       2746 = UAC71/U229/Vin (-984.5 , -81)
*       2746 = UAC71/U220/OUT (-986 , -50)
*       2752 = UAC71/U218/B (-1009.5 , -82.5)
*       2752 = UAC71/U229/Vout (-970.5 , -81)
*       2753 = UAC71/U254/Vin (-1054.5 , -125)
*       2753 = UAC71/U253/OUT (-1020 , -136.5)
*       2754 = UAC71/U253/B (-998 , -136)
*       2754 = UAC71/U246/Vout (-878.5 , -125)
*       2755 = UAC71/U218/A (-1083 , -77.5)
*       2755 = UAC71/U222/Vout (-1054 , -26.5)
*       2758 = UAC71/U245/Vout (-1104.5 , -81)
*       2758 = UAC71/U253/A (-1010.5 , -136.5)
*       2759 = UAC71/U245/Vin (-1118.5 , -81)
*       2759 = UAC71/U238/OUT (-1158 , -94)
*       2760 = UAC71/U238/B (-1145 , -82.5)
*       2760 = UAC71/U220/A (-999.5 , -38.5)
*       2760 = UAC71/C6 (-999.5 , -6.5)
*       2760 = UAC72/U254/Vout (-677 , -125)
*       2760 = UAC72/P (-676 , -152)
*       2760 = UAC71/U236/B (-874 , -82.5)
*       2760 = UAC71/C (-833.5 , -55.5)
*       2762 = UAC71/S (-1213 , -122.5)
*       2762 = r3 (-1232 , -160)
*       2762 = UAC71/U218/Vout (-1047.5 , -70.5)
*       2763 = UAC71/U254/Vout (-1040.5 , -125)
*       2763 = UAC71/P (-1039.5 , -152)



M6399 88 104 84 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
* Pins of element D6397 are shorted:
* D6397 88 88 D_lateral AREA=3.125E-016    $ (220.5 1227 220.501 1232)CMOSN6397 88 88 D_lateral AREA=3.125E-016    
M6396 88 65 2 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M6395 88 65 6 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M6394 6 1 87 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M6393 1 10 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6392 5 10 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6391 87 2 5 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M6390 84 87 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6389 88 87 86 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6388 86 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6387 94 11 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6386 88 12 11 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6385 3 65 87 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M6384 104 65 2 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6383 87 1 4 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M6382 104 10 3 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6381 1 10 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M6380 4 2 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D6378 are shorted:
* D6378 88 88 D_lateral AREA=3.125E-016    $ (206 1271.499 211 1271.5)CMOSN6378 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6377 are shorted:
* D6377 104 104 D_lateral AREA=3.125E-016    $ (137.5 1257.499 142.5 1257.5)CMOSN6377 104 104 D_lateral AREA=3.125E-016    
* Pins of element D6376 are shorted:
* D6376 88 88 D_lateral AREA=3.125E-016    $ (176 1227 176.001 1232)CMOSN6376 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6375 are shorted:
* D6375 88 88 D_lateral AREA=3.125E-016    $ (121.5 1271 121.501 1276)CMOSN6375 88 88 D_lateral AREA=3.125E-016    
M6374 88 10 8 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M6373 88 10 18 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M6372 18 7 96 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M6371 7 20 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6370 17 20 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6369 96 8 17 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M6368 11 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6367 88 94 92 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M6366 88 94 16 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M6365 91 96 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6364 16 91 244 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M6363 15 96 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6362 244 92 15 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M6361 9 10 96 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M6360 104 10 8 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6359 96 7 14 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M6358 104 20 9 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6357 7 20 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M6356 14 8 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M6355 13 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6354 13 12 11 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D6353 are shorted:
* D6353 88 88 D_lateral AREA=3.125E-016    $ (75.5 1271.499 80.5 1271.5)CMOSN6353 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6351 are shorted:
* D6351 88 88 D_lateral AREA=3.125E-016    $ (82 1227.499 87 1227.5)CMOSN6351 88 88 D_lateral AREA=3.125E-016    
M6350 88 19 20 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M6349 101 102 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6348 88 104 102 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6347 102 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6346 88 12 19 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6345 19 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6344 104 19 20 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M6343 19 12 21 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M6342 21 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D6341 are shorted:
* D6341 88 88 D_lateral AREA=3.125E-016    $ (-50.5 1227 -50.499 1232)CMOSN6341 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6340 are shorted:
* D6340 104 104 D_lateral AREA=3.125E-016    $ (7 1257.499 12 1257.5)CMOSN6340 104 104 D_lateral AREA=3.125E-016    
* Pins of element D6339 are shorted:
* D6339 88 88 D_lateral AREA=3.125E-016    $ (-50 1271 -49.999 1276)CMOSN6339 88 88 D_lateral AREA=3.125E-016    
M6338 88 65 28 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M6337 88 65 22 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M6336 22 23 27 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M6335 88 124 106 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6334 106 27 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6333 24 65 27 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M6332 104 65 28 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6331 27 23 26 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
* Pins of element D6330 are shorted:
* D6330 88 88 D_lateral AREA=3.125E-016    $ (-157.5 1271.499 -152.5 1271.5)CMOSN6330 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6329 are shorted:
* D6329 88 88 D_lateral AREA=3.125E-016    $ (-143 1227 -142.999 1232)CMOSN6329 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6328 are shorted:
* D6328 88 88 D_lateral AREA=3.125E-016    $ (-187.5 1227 -187.499 1232)CMOSN6328 88 88 D_lateral AREA=3.125E-016    
M6327 23 104 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6326 29 104 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6325 27 28 29 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M6324 88 27 110 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6323 110 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6322 35 111 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6321 31 104 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M6320 88 12 111 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6319 111 124 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6318 120 35 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M6317 23 104 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M6316 104 104 24 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6315 26 28 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M6314 104 104 31 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6313 111 12 25 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M6312 25 124 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D6311 are shorted:
* D6311 104 104 D_lateral AREA=3.125E-016    $ (-226 1257.499 -221 1257.5)CMOSN6311 104 104 D_lateral AREA=3.125E-016    
* Pins of element D6310 are shorted:
* D6310 88 88 D_lateral AREA=3.125E-016    $ (-288 1271.499 -283 1271.5)CMOSN6310 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6309 are shorted:
* D6309 88 88 D_lateral AREA=3.125E-016    $ (-242 1271 -241.999 1276)CMOSN6309 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6308 are shorted:
* D6308 88 88 D_lateral AREA=3.125E-016    $ (-281.5 1227.499 -276.5 1227.5)CMOSN6308 88 88 D_lateral AREA=3.125E-016    
M6307 88 39 40 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M6306 117 122 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6305 88 104 38 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M6304 38 30 119 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M6303 30 40 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6302 37 40 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6301 119 31 37 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M6300 88 35 36 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M6299 115 119 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6298 36 115 262 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M6297 34 119 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6296 262 120 34 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M6295 104 39 40 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M6294 32 104 119 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M6293 119 30 33 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M6292 104 40 32 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6291 30 40 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M6290 33 31 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D6289 are shorted:
* D6289 104 104 D_lateral AREA=3.125E-016    $ (-356.5 1257.499 -351.5 1257.5)CMOSN6289 104 104 D_lateral AREA=3.125E-016    
M6288 88 124 122 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6287 122 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6286 88 12 39 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6285 39 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6284 39 12 41 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M6283 41 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D6282 are shorted:
* D6282 88 88 D_lateral AREA=3.125E-016    $ (-414 1227 -413.999 1232)CMOSN6282 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6281 are shorted:
* D6281 88 88 D_lateral AREA=3.125E-016    $ (-413.5 1271 -413.499 1276)CMOSN6281 88 88 D_lateral AREA=3.125E-016    
M6280 88 65 43 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M6279 88 65 47 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M6278 47 42 128 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M6277 42 104 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6276 46 104 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6275 128 43 46 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M6274 88 148 127 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6273 127 128 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6272 88 128 126 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6271 126 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6270 44 65 128 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M6269 104 65 43 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6268 128 42 45 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M6267 104 104 44 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6266 42 104 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M6265 45 43 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D6264 are shorted:
* D6264 88 88 D_lateral AREA=3.125E-016    $ (-522 1271.499 -517 1271.5)CMOSN6264 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6263 are shorted:
* D6263 104 104 D_lateral AREA=3.125E-016    $ (-590.5 1257.499 -585.5 1257.5)CMOSN6263 104 104 D_lateral AREA=3.125E-016    
* Pins of element D6262 are shorted:
* D6262 88 88 D_lateral AREA=3.125E-016    $ (-507.5 1227 -507.499 1232)CMOSN6262 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6261 are shorted:
* D6261 88 88 D_lateral AREA=3.125E-016    $ (-552 1227 -551.999 1232)CMOSN6261 88 88 D_lateral AREA=3.125E-016    
M6260 132 136 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6259 88 104 48 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M6258 88 104 53 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M6257 53 54 143 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M6256 143 48 57 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M6255 88 12 136 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6254 136 148 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6253 88 132 131 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M6252 88 132 52 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M6251 52 140 301 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M6250 51 143 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6249 301 131 51 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M6248 55 104 143 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M6247 104 104 48 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6246 143 54 50 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M6245 50 48 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M6244 136 12 49 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M6243 49 148 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D6242 are shorted:
* D6242 88 88 D_lateral AREA=3.125E-016    $ (-652.5 1271.499 -647.5 1271.5)CMOSN6242 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6241 are shorted:
* D6241 88 88 D_lateral AREA=3.125E-016    $ (-606.5 1271 -606.499 1276)CMOSN6241 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6240 are shorted:
* D6240 88 88 D_lateral AREA=3.125E-016    $ (-646 1227.499 -641 1227.5)CMOSN6240 88 88 D_lateral AREA=3.125E-016    
M6239 88 58 56 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M6238 142 144 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6237 88 148 144 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6236 54 56 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6235 57 56 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6234 88 12 58 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6233 140 143 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6232 104 58 56 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M6231 54 56 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M6230 104 56 55 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D6228 are shorted:
* D6228 88 88 D_lateral AREA=3.125E-016    $ (-778.5 1227 -778.499 1232)CMOSN6228 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6227 are shorted:
* D6227 104 104 D_lateral AREA=3.125E-016    $ (-721 1257.499 -716 1257.5)CMOSN6227 104 104 D_lateral AREA=3.125E-016    
* Pins of element D6226 are shorted:
* D6226 88 88 D_lateral AREA=3.125E-016    $ (-778 1271 -777.999 1276)CMOSN6226 88 88 D_lateral AREA=3.125E-016    
M6225 144 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6224 58 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6223 60 65 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M6222 88 71 146 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6221 146 152 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6220 59 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6219 59 12 58 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6218 104 65 60 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D6217 are shorted:
* D6217 88 88 D_lateral AREA=3.125E-016    $ (-885.5 1271.499 -880.5 1271.5)CMOSN6217 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6216 are shorted:
* D6216 88 88 D_lateral AREA=3.125E-016    $ (-871 1227 -870.999 1232)CMOSN6216 88 88 D_lateral AREA=3.125E-016    
M6215 88 65 67 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M6214 67 61 152 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M6213 61 104 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6212 66 104 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6211 152 60 66 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M6210 88 152 151 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6209 151 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6208 159 153 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6207 88 12 153 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6206 153 71 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6205 62 65 152 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M6204 152 61 64 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M6203 104 104 62 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6202 61 104 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M6201 64 60 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M6200 153 12 63 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M6199 63 71 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D6198 are shorted:
* D6198 104 104 D_lateral AREA=3.125E-016    $ (-954 1257.499 -949 1257.5)CMOSN6198 104 104 D_lateral AREA=3.125E-016    
* Pins of element D6197 are shorted:
* D6197 88 88 D_lateral AREA=3.125E-016    $ (-915.5 1227 -915.499 1232)CMOSN6197 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6196 are shorted:
* D6196 88 88 D_lateral AREA=3.125E-016    $ (-970 1271 -969.999 1276)CMOSN6196 88 88 D_lateral AREA=3.125E-016    
M6195 88 104 69 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M6194 88 104 76 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M6193 76 68 162 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M6192 68 78 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6191 75 78 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6190 162 69 75 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M6189 88 159 157 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M6188 88 159 74 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M6187 156 162 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6186 74 156 337 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M6185 73 162 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6184 337 157 73 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M6183 70 104 162 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M6182 104 104 69 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6181 162 68 72 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M6180 104 78 70 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6179 68 78 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M6178 72 69 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D6177 are shorted:
* D6177 88 88 D_lateral AREA=3.125E-016    $ (-1016 1271.499 -1011 1271.5)CMOSN6177 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6176 are shorted:
* D6176 104 104 D_lateral AREA=3.125E-016    $ (-1084.5 1257.499 -1079.5 1257.5)CMOSN6176 104 104 D_lateral AREA=3.125E-016    
* Pins of element D6175 are shorted:
* D6175 88 88 D_lateral AREA=3.125E-016    $ (-1009.5 1227.499 -1004.5 1227.5)CMOSN6175 88 88 D_lateral AREA=3.125E-016    
M6174 88 77 78 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M6173 165 166 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6172 88 71 166 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6171 166 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6170 88 12 77 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6169 77 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6168 104 77 78 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M6167 77 12 79 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M6166 79 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D6165 are shorted:
* D6165 88 88 D_lateral AREA=3.125E-016    $ (-1142 1227 -1141.999 1232)CMOSN6165 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6164 are shorted:
* D6164 88 88 D_lateral AREA=3.125E-016    $ (-1141.5 1271 -1141.499 1276)CMOSN6164 88 88 D_lateral AREA=3.125E-016    
M6162 88 88 172 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6161 172 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6160 12 80 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M6159 81 491 88 88 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M6158 80 174 81 88 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M6156 12 80 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6155 80 491 104 104 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M6154 104 174 80 104 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
* Pins of element D6153 are shorted:
* D6153 88 88 D_lateral AREA=3.125E-016    $ (-1414 1225.5 -1413.999 1230.5)CMOSN6153 88 88 D_lateral AREA=3.125E-016    
M6152 88 183 181 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6151 181 182 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6149 10 82 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M6148 88 183 82 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M6147 82 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6146 10 82 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6145 82 183 83 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M6144 83 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D6143 are shorted:
* D6143 88 88 D_lateral AREA=3.125E-016    $ (-1498 1225.5 -1497.999 1230.5)CMOSN6143 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6142 are shorted:
* D6142 88 88 D_lateral AREA=3.125E-016    $ (-1527 1271 -1526.999 1276)CMOSN6142 88 88 D_lateral AREA=3.125E-016    
M6141 95 84 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6140 95 84 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M6138 88 85 99 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M6137 85 86 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6136 104 85 98 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M6135 85 86 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M6134 90 87 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6133 90 104 84 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6132 86 87 89 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M6131 89 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6130 94 11 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D6129 are shorted:
* D6129 88 88 D_lateral AREA=3.125E-016    $ (126.5 1182 126.501 1187)CMOSN6129 88 88 D_lateral AREA=3.125E-016    
* Pins of element D6128 are shorted:
* D6128 104 104 D_lateral AREA=3.125E-016    $ (127.999 1165 128 1170)CMOSN6128 104 104 D_lateral AREA=3.125E-016    
M6127 124 98 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6126 99 95 100 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M6125 100 101 98 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M6124 124 98 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M6123 98 95 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M6122 104 101 98 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M6121 93 94 244 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M6120 104 94 92 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6119 244 91 97 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M6118 104 96 93 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6117 91 96 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M6116 97 92 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D6115 are shorted:
* D6115 104 104 D_lateral AREA=3.125E-016    $ (13.5 1213.499 18.5 1213.5)CMOSN6115 104 104 D_lateral AREA=3.125E-016    
M6114 101 102 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M6113 102 104 105 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M6112 105 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6111 108 106 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6110 108 106 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M6109 106 124 107 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M6108 107 27 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6107 113 108 114 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M6106 88 109 113 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M6105 114 117 118 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M6104 109 110 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6103 118 108 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M6102 104 109 118 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M6101 104 117 118 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M6100 109 110 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M6099 110 27 112 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M6098 112 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6097 35 111 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M6096 104 35 120 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D6095 are shorted:
* D6095 104 104 D_lateral AREA=3.125E-016    $ (-235.501 1165 -235.5 1170)CMOSN6095 104 104 D_lateral AREA=3.125E-016    
* Pins of element D6094 are shorted:
* D6094 88 88 D_lateral AREA=3.125E-016    $ (-237 1182 -236.999 1187)CMOSN6094 88 88 D_lateral AREA=3.125E-016    
M6093 148 118 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6092 148 118 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M6091 117 122 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M6090 116 35 262 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M6089 262 115 121 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M6088 104 119 116 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6087 115 119 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M6086 121 120 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D6085 are shorted:
* D6085 104 104 D_lateral AREA=3.125E-016    $ (-350 1213.499 -345 1213.5)CMOSN6085 104 104 D_lateral AREA=3.125E-016    
M6084 122 124 125 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M6083 125 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6082 135 126 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6081 134 127 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6080 135 126 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M6079 134 127 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M6078 127 148 130 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M6077 130 128 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6076 126 128 129 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M6075 129 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6074 71 133 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6073 138 134 139 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M6072 88 135 138 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M6071 139 142 133 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M6070 71 133 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M6069 133 134 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M6068 104 135 133 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M6067 104 142 133 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M6066 132 136 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M6065 141 132 301 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M6064 104 132 131 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6063 301 140 137 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M6061 137 131 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D6060 are shorted:
* D6060 104 104 D_lateral AREA=3.125E-016    $ (-600.001 1165 -600 1170)CMOSN6060 104 104 D_lateral AREA=3.125E-016    
* Pins of element D6059 are shorted:
* D6059 88 88 D_lateral AREA=3.125E-016    $ (-601.5 1182 -601.499 1187)CMOSN6059 88 88 D_lateral AREA=3.125E-016    
M6058 142 144 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M6056 140 143 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M6055 141 143 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
* Pins of element D6054 are shorted:
* D6054 104 104 D_lateral AREA=3.125E-016    $ (-714.5 1213.499 -709.5 1213.5)CMOSN6054 104 104 D_lateral AREA=3.125E-016    
M6053 161 146 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6052 149 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6051 149 148 144 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6050 161 146 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M6049 146 71 147 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M6048 147 152 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6047 155 161 164 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M6046 88 150 155 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M6045 150 151 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6044 160 161 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M6043 104 150 160 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M6042 150 151 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M6041 151 152 154 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M6040 154 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6039 159 153 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D6038 are shorted:
* D6038 104 104 D_lateral AREA=3.125E-016    $ (-963.501 1165 -963.5 1170)CMOSN6038 104 104 D_lateral AREA=3.125E-016    
* Pins of element D6037 are shorted:
* D6037 88 88 D_lateral AREA=3.125E-016    $ (-965 1182 -964.999 1187)CMOSN6037 88 88 D_lateral AREA=3.125E-016    
M6036 179 160 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M6035 164 165 160 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M6034 179 160 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M6033 104 165 160 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M6032 158 159 337 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M6031 104 159 157 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6030 337 156 163 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M6029 104 162 158 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6028 156 162 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M6027 163 157 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D6026 are shorted:
* D6026 104 104 D_lateral AREA=3.125E-016    $ (-1078 1213.499 -1073 1213.5)CMOSN6026 104 104 D_lateral AREA=3.125E-016    
M6025 165 166 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M6024 166 71 168 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M6023 168 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6022 65 172 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M6020 65 172 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D6019 are shorted:
* D6019 88 88 D_lateral AREA=3.125E-016    $ (-1391 1180.999 -1386 1181)CMOSN6019 88 88 D_lateral AREA=3.125E-016    
M6018 88 65 170 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M6017 88 65 178 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M6016 178 169 186 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M6015 169 173 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6014 177 173 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6013 186 170 177 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M6011 174 181 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M6010 171 65 186 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M6009 170 65 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M6008 186 169 176 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M6007 104 173 171 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6006 169 173 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M6005 176 170 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M6003 172 88 175 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M6002 175 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M6001 174 181 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D6000 are shorted:
* D6000 104 104 D_lateral AREA=3.125E-016    $ (-1459.5 1166.999 -1454.5 1167)CMOSN6000 104 104 D_lateral AREA=3.125E-016    
M5999 88 180 173 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M5998 88 179 180 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5997 180 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5996 182 491 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M5995 104 180 173 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5994 180 179 185 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5993 185 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5992 181 183 184 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5991 184 182 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5990 182 491 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D5989 are shorted:
* D5989 88 88 D_lateral AREA=3.125E-016    $ (-1519 1180.5 -1518.999 1185.5)CMOSN5989 88 88 D_lateral AREA=3.125E-016    
M5987 88 104 363 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
* Pins of element D5984 are shorted:
* D5984 88 88 D_lateral AREA=3.125E-016    $ (220 1064.5 220.001 1069.5)CMOSN5984 88 88 D_lateral AREA=3.125E-016    
M5983 88 469 188 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5982 88 469 195 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5981 195 187 190 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5980 187 353 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5979 194 353 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5978 190 188 194 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5976 363 190 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5975 88 190 365 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5974 365 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5973 202 204 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5972 88 206 204 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5971 189 469 190 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5970 104 469 188 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5969 190 187 193 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5968 104 353 189 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5967 187 353 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5966 193 188 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M5965 192 190 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5964 192 104 363 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5963 365 190 191 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5962 191 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5961 202 204 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D5959 are shorted:
* D5959 88 88 D_lateral AREA=3.125E-016    $ (205.5 1108.999 210.5 1109)CMOSN5959 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5958 are shorted:
* D5958 104 104 D_lateral AREA=3.125E-016    $ (137 1094.999 142 1095)CMOSN5958 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5957 are shorted:
* D5957 88 88 D_lateral AREA=3.125E-016    $ (175.5 1064.5 175.501 1069.5)CMOSN5957 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5956 are shorted:
* D5956 88 88 D_lateral AREA=3.125E-016    $ (121 1108.5 121.001 1113.5)CMOSN5956 88 88 D_lateral AREA=3.125E-016    
M5954 88 353 197 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5953 88 353 212 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5952 212 196 203 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5951 196 214 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5950 211 214 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5949 203 197 211 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5948 204 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5947 88 202 200 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5946 88 202 210 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5945 210 199 400 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5944 199 203 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5943 209 203 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5942 400 200 209 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5941 198 353 203 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5940 104 353 197 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5939 203 196 208 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5938 104 214 198 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5937 196 214 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5936 208 197 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M5935 207 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5934 207 206 204 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5933 201 202 400 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5932 104 202 200 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5931 400 199 205 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5930 104 203 201 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5929 199 203 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5928 205 200 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D5927 are shorted:
* D5927 88 88 D_lateral AREA=3.125E-016    $ (75 1108.999 80 1109)CMOSN5927 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5925 are shorted:
* D5925 88 88 D_lateral AREA=3.125E-016    $ (81.5 1064.999 86.5 1065)CMOSN5925 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5924 are shorted:
* D5924 104 104 D_lateral AREA=3.125E-016    $ (13 1050.999 18 1051)CMOSN5924 104 104 D_lateral AREA=3.125E-016    
M5923 88 213 214 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M5922 215 216 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5921 88 104 216 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5920 216 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5919 88 206 213 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5918 213 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5917 104 213 214 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M5916 215 216 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5915 216 104 218 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5914 218 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5913 213 206 217 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5912 217 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5911 are shorted:
* D5911 88 88 D_lateral AREA=3.125E-016    $ (-51 1064.5 -50.999 1069.5)CMOSN5911 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5910 are shorted:
* D5910 104 104 D_lateral AREA=3.125E-016    $ (6.5 1094.999 11.5 1095)CMOSN5910 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5909 are shorted:
* D5909 88 88 D_lateral AREA=3.125E-016    $ (-50.5 1108.5 -50.499 1113.5)CMOSN5909 88 88 D_lateral AREA=3.125E-016    
M5908 88 469 228 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5907 88 469 220 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5906 220 221 227 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5904 88 247 380 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5903 380 227 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5902 222 469 227 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5901 104 469 228 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5900 227 221 226 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5899 380 247 219 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5898 219 227 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5897 are shorted:
* D5897 88 88 D_lateral AREA=3.125E-016    $ (-158 1108.999 -153 1109)CMOSN5897 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5896 are shorted:
* D5896 88 88 D_lateral AREA=3.125E-016    $ (-143.5 1064.5 -143.499 1069.5)CMOSN5896 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5895 are shorted:
* D5895 88 88 D_lateral AREA=3.125E-016    $ (-188 1064.5 -187.999 1069.5)CMOSN5895 88 88 D_lateral AREA=3.125E-016    
M5894 221 244 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5893 229 244 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5892 227 228 229 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5890 88 227 386 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5889 386 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5888 238 223 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5886 88 206 223 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5885 223 247 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5884 236 238 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M5883 221 244 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5882 104 244 222 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5881 226 228 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M5880 386 227 225 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5879 225 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5878 238 223 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5877 104 244 231 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5876 223 206 224 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5875 224 247 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5874 104 238 236 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D5873 are shorted:
* D5873 104 104 D_lateral AREA=3.125E-016    $ (-226.5 1094.999 -221.5 1095)CMOSN5873 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5872 are shorted:
* D5872 88 88 D_lateral AREA=3.125E-016    $ (-288.5 1108.999 -283.5 1109)CMOSN5872 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5871 are shorted:
* D5871 88 88 D_lateral AREA=3.125E-016    $ (-242.5 1108.5 -242.499 1113.5)CMOSN5871 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5870 are shorted:
* D5870 88 88 D_lateral AREA=3.125E-016    $ (-282 1064.999 -277 1065)CMOSN5870 88 88 D_lateral AREA=3.125E-016    
M5869 88 245 246 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M5867 395 248 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5866 231 244 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M5865 88 244 243 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5864 243 230 235 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5863 230 246 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5862 242 246 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5861 235 231 242 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5860 88 238 241 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5859 241 233 558 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5858 233 235 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5857 240 235 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5856 558 236 240 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5855 104 245 246 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M5854 395 248 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5853 232 244 235 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5852 235 230 239 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5851 104 246 232 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5850 230 246 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5849 239 231 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M5848 234 238 558 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5847 558 233 237 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5846 104 235 234 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5845 233 235 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5844 237 236 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D5843 are shorted:
* D5843 104 104 D_lateral AREA=3.125E-016    $ (-357 1094.999 -352 1095)CMOSN5843 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5842 are shorted:
* D5842 104 104 D_lateral AREA=3.125E-016    $ (-350.5 1050.999 -345.5 1051)CMOSN5842 104 104 D_lateral AREA=3.125E-016    
M5841 88 247 248 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5840 248 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5839 88 206 245 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5838 245 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5837 248 247 250 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5836 250 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5835 245 206 249 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5834 249 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5833 are shorted:
* D5833 88 88 D_lateral AREA=3.125E-016    $ (-414.5 1064.5 -414.499 1069.5)CMOSN5833 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5832 are shorted:
* D5832 88 88 D_lateral AREA=3.125E-016    $ (-414 1108.5 -413.999 1113.5)CMOSN5832 88 88 D_lateral AREA=3.125E-016    
M5831 88 469 252 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5830 88 469 259 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5829 259 251 254 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5828 251 262 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5827 258 262 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5826 254 252 258 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5823 88 282 405 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5822 405 254 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5821 88 254 404 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5820 404 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5819 253 469 254 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5818 104 469 252 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5817 254 251 257 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5816 104 262 253 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5815 251 262 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5814 257 252 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M5813 405 282 256 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5812 256 254 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5811 404 254 255 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5810 255 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5809 are shorted:
* D5809 88 88 D_lateral AREA=3.125E-016    $ (-522.5 1108.999 -517.5 1109)CMOSN5809 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5808 are shorted:
* D5808 104 104 D_lateral AREA=3.125E-016    $ (-591 1094.999 -586 1095)CMOSN5808 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5807 are shorted:
* D5807 88 88 D_lateral AREA=3.125E-016    $ (-508 1064.5 -507.999 1069.5)CMOSN5807 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5806 are shorted:
* D5806 88 88 D_lateral AREA=3.125E-016    $ (-552.5 1064.5 -552.499 1069.5)CMOSN5806 88 88 D_lateral AREA=3.125E-016    
M5804 263 264 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5803 88 262 260 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5802 88 262 270 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5801 270 271 276 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5800 276 260 277 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5799 88 206 264 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5798 264 282 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5797 88 263 261 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5796 88 263 269 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5795 269 273 589 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5794 268 276 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5793 589 261 268 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5792 263 264 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5791 272 262 276 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5790 104 262 260 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5789 276 271 267 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5788 267 260 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M5787 264 206 266 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5786 266 282 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5785 274 263 589 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5784 104 263 261 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5783 589 273 265 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5781 265 261 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D5780 are shorted:
* D5780 88 88 D_lateral AREA=3.125E-016    $ (-653 1108.999 -648 1109)CMOSN5780 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5779 are shorted:
* D5779 88 88 D_lateral AREA=3.125E-016    $ (-607 1108.5 -606.999 1113.5)CMOSN5779 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5778 are shorted:
* D5778 88 88 D_lateral AREA=3.125E-016    $ (-646.5 1064.999 -641.5 1065)CMOSN5778 88 88 D_lateral AREA=3.125E-016    
M5777 88 278 275 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M5776 419 279 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5775 88 282 279 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5774 271 275 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5773 277 275 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5772 88 206 278 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5771 273 276 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5770 104 278 275 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M5769 419 279 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5767 271 275 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5766 104 275 272 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5764 273 276 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5763 274 276 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
* Pins of element D5762 are shorted:
* D5762 88 88 D_lateral AREA=3.125E-016    $ (-779 1064.5 -778.999 1069.5)CMOSN5762 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5761 are shorted:
* D5761 104 104 D_lateral AREA=3.125E-016    $ (-721.5 1094.999 -716.5 1095)CMOSN5761 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5760 are shorted:
* D5760 88 88 D_lateral AREA=3.125E-016    $ (-778.5 1108.5 -778.499 1113.5)CMOSN5760 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5759 are shorted:
* D5759 104 104 D_lateral AREA=3.125E-016    $ (-715 1050.999 -710 1051)CMOSN5759 104 104 D_lateral AREA=3.125E-016    
M5758 279 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5757 278 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5756 284 469 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M5754 88 300 422 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5753 422 287 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5752 283 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5751 283 282 279 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5750 281 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5749 281 206 278 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5748 104 469 284 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5747 422 300 280 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5746 280 287 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5745 are shorted:
* D5745 88 88 D_lateral AREA=3.125E-016    $ (-886 1108.999 -881 1109)CMOSN5745 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5744 are shorted:
* D5744 88 88 D_lateral AREA=3.125E-016    $ (-871.5 1064.5 -871.499 1069.5)CMOSN5744 88 88 D_lateral AREA=3.125E-016    
M5743 88 469 293 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5742 293 285 287 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5741 285 301 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5740 292 301 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5739 287 284 292 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5737 88 287 427 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5736 427 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5735 302 288 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5734 88 206 288 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5733 288 300 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5732 286 469 287 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5731 287 285 291 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5730 104 301 286 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5729 285 301 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5728 291 284 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M5727 427 287 290 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5726 290 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5725 302 288 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5724 288 206 289 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5723 289 300 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5722 are shorted:
* D5722 104 104 D_lateral AREA=3.125E-016    $ (-954.5 1094.999 -949.5 1095)CMOSN5722 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5721 are shorted:
* D5721 88 88 D_lateral AREA=3.125E-016    $ (-916 1064.5 -915.999 1069.5)CMOSN5721 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5720 are shorted:
* D5720 88 88 D_lateral AREA=3.125E-016    $ (-970.5 1108.5 -970.499 1113.5)CMOSN5720 88 88 D_lateral AREA=3.125E-016    
M5718 88 301 295 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5717 88 301 309 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5716 309 294 303 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5715 294 311 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5714 308 311 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5713 303 295 308 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5712 88 302 298 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5711 88 302 307 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5710 307 297 460 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5709 297 303 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5708 306 303 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5707 460 298 306 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5706 296 301 303 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5705 104 301 295 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5704 303 294 305 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5703 104 311 296 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5702 294 311 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5701 305 295 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M5700 299 302 460 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5699 104 302 298 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5698 460 297 304 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5697 104 303 299 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5696 297 303 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5695 304 298 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D5694 are shorted:
* D5694 88 88 D_lateral AREA=3.125E-016    $ (-1016.5 1108.999 -1011.5 1109)CMOSN5694 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5693 are shorted:
* D5693 104 104 D_lateral AREA=3.125E-016    $ (-1085 1094.999 -1080 1095)CMOSN5693 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5692 are shorted:
* D5692 88 88 D_lateral AREA=3.125E-016    $ (-1010 1064.999 -1005 1065)CMOSN5692 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5691 are shorted:
* D5691 104 104 D_lateral AREA=3.125E-016    $ (-1078.5 1050.999 -1073.5 1051)CMOSN5691 104 104 D_lateral AREA=3.125E-016    
M5690 88 310 311 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M5689 312 313 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5688 88 300 313 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5687 313 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5686 88 206 310 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5685 310 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5684 104 310 311 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M5683 312 313 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5682 313 300 315 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5681 315 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5680 310 206 314 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5679 314 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5678 are shorted:
* D5678 88 88 D_lateral AREA=3.125E-016    $ (-1142.5 1064.5 -1142.499 1069.5)CMOSN5678 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5677 are shorted:
* D5677 88 88 D_lateral AREA=3.125E-016    $ (-1142 1108.5 -1141.999 1113.5)CMOSN5677 88 88 D_lateral AREA=3.125E-016    
M5676 88 469 316 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5675 88 469 320 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5674 320 321 325 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5672 325 316 319 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5670 88 345 443 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5669 443 325 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5668 88 325 451 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5667 322 469 325 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5666 104 469 316 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5665 325 321 318 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5664 318 316 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M5663 443 345 317 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5662 317 325 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5660 are shorted:
* D5660 88 88 D_lateral AREA=3.125E-016    $ (-1250 1108.999 -1245 1109)CMOSN5660 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5659 are shorted:
* D5659 88 88 D_lateral AREA=3.125E-016    $ (-1235.5 1064.5 -1235.499 1069.5)CMOSN5659 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5658 are shorted:
* D5658 88 88 D_lateral AREA=3.125E-016    $ (-1280 1064.5 -1279.999 1069.5)CMOSN5658 88 88 D_lateral AREA=3.125E-016    
M5657 321 337 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5656 88 337 319 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5654 451 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5653 335 323 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5652 341 337 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M5651 88 206 323 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5650 323 345 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5649 338 335 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M5648 321 337 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5647 104 337 322 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5646 326 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5645 326 325 451 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5644 335 323 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5643 104 337 341 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5642 323 206 324 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5641 324 345 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5639 104 335 338 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D5638 are shorted:
* D5638 104 104 D_lateral AREA=3.125E-016    $ (-1318.5 1094.999 -1313.5 1095)CMOSN5638 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5637 are shorted:
* D5637 88 88 D_lateral AREA=3.125E-016    $ (-1380.5 1108.999 -1375.5 1109)CMOSN5637 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5636 are shorted:
* D5636 88 88 D_lateral AREA=3.125E-016    $ (-1334.5 1108.5 -1334.499 1113.5)CMOSN5636 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5635 are shorted:
* D5635 88 88 D_lateral AREA=3.125E-016    $ (-1374 1064.999 -1369 1065)CMOSN5635 88 88 D_lateral AREA=3.125E-016    
M5634 88 344 331 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M5632 457 346 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5631 88 337 343 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5630 343 327 332 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5629 327 331 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5628 342 331 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5627 332 341 342 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5626 88 335 340 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5625 340 329 333 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5624 329 332 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5623 339 332 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5622 333 338 339 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5621 104 344 331 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M5620 457 346 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5619 328 337 332 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5618 332 327 336 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5617 104 331 328 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5616 327 331 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5615 336 341 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M5614 333 335 330 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=1.75p PS=5.5u    
M5613 333 329 334 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5612 104 332 330 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5611 329 332 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5610 334 338 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D5609 are shorted:
* D5609 104 104 D_lateral AREA=3.125E-016    $ (-1449 1094.999 -1444 1095)CMOSN5609 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5608 are shorted:
* D5608 104 104 D_lateral AREA=3.125E-016    $ (-1442.5 1050.999 -1437.5 1051)CMOSN5608 104 104 D_lateral AREA=3.125E-016    
M5607 88 345 346 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5606 346 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5605 88 206 344 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5604 344 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5603 346 345 348 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5602 348 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5601 344 206 347 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5600 347 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5599 are shorted:
* D5599 88 88 D_lateral AREA=3.125E-016    $ (-1506.5 1064.5 -1506.499 1069.5)CMOSN5599 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5598 are shorted:
* D5598 88 88 D_lateral AREA=3.125E-016    $ (-1506 1108.5 -1505.999 1113.5)CMOSN5598 88 88 D_lateral AREA=3.125E-016    
M5597 469 349 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M5596 88 186 349 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5595 206 352 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M5594 469 349 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5592 206 352 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D5591 are shorted:
* D5591 88 88 D_lateral AREA=3.125E-016    $ (-1779.5 1063 -1779.499 1068)CMOSN5591 88 88 D_lateral AREA=3.125E-016    
M5590 349 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5589 356 491 88 88 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M5588 352 351 356 88 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M5587 351 350 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M5586 88 357 350 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5585 350 359 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5584 353 358 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M5583 355 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5582 355 186 349 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5581 352 491 104 104 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M5580 104 351 352 104 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M5579 351 350 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5578 350 357 354 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5577 354 359 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5576 353 358 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D5575 are shorted:
* D5575 88 88 D_lateral AREA=3.125E-016    $ (-1863.5 1063 -1863.499 1068)CMOSN5575 88 88 D_lateral AREA=3.125E-016    
M5574 359 491 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M5573 88 357 358 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5572 358 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5571 359 491 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5570 358 357 360 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5569 360 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5568 are shorted:
* D5568 88 88 D_lateral AREA=3.125E-016    $ (-1892.5 1108.5 -1892.499 1113.5)CMOSN5568 88 88 D_lateral AREA=3.125E-016    
M5567 371 363 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5566 371 363 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5564 88 430 492 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5563 88 430 368 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5562 368 361 494 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5561 361 506 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5560 367 506 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5559 494 492 367 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5558 88 503 508 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5557 88 364 375 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M5556 364 365 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5555 362 430 494 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5554 104 430 492 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5553 494 361 366 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5552 104 506 362 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5551 361 506 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5550 366 492 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M5548 104 364 372 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M5547 364 365 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D5546 are shorted:
* D5546 88 88 D_lateral AREA=3.125E-016    $ (205 946.499 210 946.5)CMOSN5546 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5545 are shorted:
* D5545 104 104 D_lateral AREA=3.125E-016    $ (136.5 932.499 141.5 932.5)CMOSN5545 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5544 are shorted:
* D5544 88 88 D_lateral AREA=3.125E-016    $ (120.5 946 120.501 951)CMOSN5544 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5543 are shorted:
* D5543 88 88 D_lateral AREA=3.125E-016    $ (126 1019.5 126.001 1024.5)CMOSN5543 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5542 are shorted:
* D5542 104 104 D_lateral AREA=3.125E-016    $ (127.499 1002.5 127.5 1007.5)CMOSN5542 104 104 D_lateral AREA=3.125E-016    
M5541 88 506 502 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5540 88 506 378 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5539 378 369 507 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5538 369 518 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5537 377 518 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5536 507 502 377 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5535 508 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5534 247 372 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5533 375 371 376 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M5532 376 215 372 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M5531 370 506 507 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5530 104 506 502 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5529 507 369 374 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5528 104 518 370 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5527 369 518 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5526 374 502 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M5525 373 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5524 373 503 508 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5523 247 372 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5522 372 371 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M5521 104 215 372 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
* Pins of element D5520 are shorted:
* D5520 88 88 D_lateral AREA=3.125E-016    $ (74.5 946.499 79.5 946.5)CMOSN5520 88 88 D_lateral AREA=3.125E-016    
M5518 88 515 518 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M5517 88 503 515 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5516 515 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5515 104 515 518 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M5514 515 503 379 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5513 379 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5512 are shorted:
* D5512 104 104 D_lateral AREA=3.125E-016    $ (6 932.499 11 932.5)CMOSN5512 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5511 are shorted:
* D5511 88 88 D_lateral AREA=3.125E-016    $ (-51 946 -50.999 951)CMOSN5511 88 88 D_lateral AREA=3.125E-016    
M5510 88 430 522 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5509 88 430 381 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5508 381 382 391 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5507 384 380 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5506 383 430 391 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5505 104 430 522 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5504 391 382 388 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5503 384 380 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D5502 are shorted:
* D5502 88 88 D_lateral AREA=3.125E-016    $ (-158.5 946.499 -153.5 946.5)CMOSN5502 88 88 D_lateral AREA=3.125E-016    
M5501 382 400 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5500 392 400 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5499 391 522 392 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5497 88 503 526 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5496 526 543 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5495 389 384 390 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M5494 88 385 389 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M5493 390 395 396 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M5492 385 386 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5491 382 400 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5490 104 400 383 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5489 388 522 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M5488 104 400 532 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5487 526 503 387 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5486 387 543 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5485 396 384 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M5484 104 385 396 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M5483 104 395 396 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M5482 385 386 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D5481 are shorted:
* D5481 104 104 D_lateral AREA=3.125E-016    $ (-227 932.499 -222 932.5)CMOSN5481 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5480 are shorted:
* D5480 88 88 D_lateral AREA=3.125E-016    $ (-289 946.499 -284 946.5)CMOSN5480 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5479 are shorted:
* D5479 88 88 D_lateral AREA=3.125E-016    $ (-243 946 -242.999 951)CMOSN5479 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5478 are shorted:
* D5478 104 104 D_lateral AREA=3.125E-016    $ (-236.001 1002.5 -236 1007.5)CMOSN5478 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5477 are shorted:
* D5477 88 88 D_lateral AREA=3.125E-016    $ (-237.5 1019.5 -237.499 1024.5)CMOSN5477 88 88 D_lateral AREA=3.125E-016    
M5476 88 544 542 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M5475 532 400 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M5474 88 400 399 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5473 399 393 535 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5472 393 542 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5471 398 542 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5470 535 532 398 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5469 282 396 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5468 104 544 542 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M5467 394 400 535 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5466 535 393 397 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5465 104 542 394 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5464 393 542 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5463 397 532 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M5462 282 396 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D5461 are shorted:
* D5461 104 104 D_lateral AREA=3.125E-016    $ (-357.5 932.499 -352.5 932.5)CMOSN5461 104 104 D_lateral AREA=3.125E-016    
M5460 88 503 544 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5459 544 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5458 544 503 401 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5457 401 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5456 are shorted:
* D5456 88 88 D_lateral AREA=3.125E-016    $ (-414.5 946 -414.499 951)CMOSN5456 88 88 D_lateral AREA=3.125E-016    
M5455 411 404 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5454 410 405 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5453 88 430 546 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5452 88 430 408 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5451 408 402 547 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5450 402 558 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5449 407 558 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5448 547 546 407 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5447 411 404 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5446 410 405 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5445 403 430 547 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5444 104 430 546 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5443 547 402 406 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5442 104 558 403 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5441 402 558 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5440 406 546 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D5439 are shorted:
* D5439 88 88 D_lateral AREA=3.125E-016    $ (-523 946.499 -518 946.5)CMOSN5439 88 88 D_lateral AREA=3.125E-016    
M5437 300 409 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5436 415 410 416 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M5435 88 411 415 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M5434 416 419 409 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M5433 88 558 420 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5432 88 558 414 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5431 414 417 569 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5429 88 503 557 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5428 557 573 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5427 300 409 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5426 409 410 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M5425 104 411 409 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M5424 104 419 409 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M5423 418 558 569 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5422 104 558 420 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5421 569 417 413 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5420 104 420 413 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=187.5f PS=1.25u    
M5419 557 503 412 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5418 412 573 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5417 are shorted:
* D5417 104 104 D_lateral AREA=3.125E-016    $ (-600.501 1002.5 -600.5 1007.5)CMOSN5417 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5416 are shorted:
* D5416 88 88 D_lateral AREA=3.125E-016    $ (-602 1019.5 -601.999 1024.5)CMOSN5416 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5415 are shorted:
* D5415 104 104 D_lateral AREA=3.125E-016    $ (-591.5 932.499 -586.5 932.5)CMOSN5415 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5414 are shorted:
* D5414 88 88 D_lateral AREA=3.125E-016    $ (-653.5 946.499 -648.5 946.5)CMOSN5414 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5413 are shorted:
* D5413 88 88 D_lateral AREA=3.125E-016    $ (-607.5 946 -607.499 951)CMOSN5413 88 88 D_lateral AREA=3.125E-016    
M5412 88 566 568 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M5411 417 568 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5410 421 568 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5409 421 420 569 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5408 88 503 566 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5407 104 566 568 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M5406 417 568 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5405 104 568 418 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D5403 are shorted:
* D5403 104 104 D_lateral AREA=3.125E-016    $ (-722 932.499 -717 932.5)CMOSN5403 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5402 are shorted:
* D5402 88 88 D_lateral AREA=3.125E-016    $ (-779 946 -778.999 951)CMOSN5402 88 88 D_lateral AREA=3.125E-016    
M5401 566 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5400 575 430 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M5399 437 422 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5398 423 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5397 423 503 566 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5396 104 430 575 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5395 437 422 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D5394 are shorted:
* D5394 88 88 D_lateral AREA=3.125E-016    $ (-886.5 946.499 -881.5 946.5)CMOSN5394 88 88 D_lateral AREA=3.125E-016    
M5393 88 430 433 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5392 433 424 577 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5391 424 589 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5390 432 589 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5389 577 575 432 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5388 88 503 579 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5387 579 599 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5386 431 437 439 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M5385 88 426 431 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M5384 426 427 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5383 425 430 577 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5382 577 424 429 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5381 104 589 425 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5380 424 589 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5379 429 575 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M5378 579 503 428 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5377 104 599 428 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5376 436 437 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M5375 104 426 436 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M5374 426 427 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D5373 are shorted:
* D5373 104 104 D_lateral AREA=3.125E-016    $ (-955 932.499 -950 932.5)CMOSN5373 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5372 are shorted:
* D5372 88 88 D_lateral AREA=3.125E-016    $ (-971 946 -970.999 951)CMOSN5372 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5371 are shorted:
* D5371 88 88 D_lateral AREA=3.125E-016    $ (-965.5 1019.5 -965.499 1024.5)CMOSN5371 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5370 are shorted:
* D5370 104 104 D_lateral AREA=3.125E-016    $ (-964.001 1002.5 -964 1007.5)CMOSN5370 104 104 D_lateral AREA=3.125E-016    
M5369 88 589 585 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5368 88 589 441 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5367 441 434 590 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5366 434 598 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5365 440 598 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5364 590 585 440 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5363 345 436 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5362 439 312 436 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M5361 435 589 590 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5360 104 589 585 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5359 590 434 438 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5358 104 598 435 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5357 434 598 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5356 438 585 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M5355 345 436 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5354 104 312 436 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
* Pins of element D5353 are shorted:
* D5353 88 88 D_lateral AREA=3.125E-016    $ (-1017 946.499 -1012 946.5)CMOSN5353 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5352 are shorted:
* D5352 104 104 D_lateral AREA=3.125E-016    $ (-1085.5 932.499 -1080.5 932.5)CMOSN5352 104 104 D_lateral AREA=3.125E-016    
M5351 88 595 598 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M5350 88 503 595 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5349 595 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5348 104 595 598 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M5347 595 503 442 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5346 442 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5345 are shorted:
* D5345 88 88 D_lateral AREA=3.125E-016    $ (-1142.5 946 -1142.499 951)CMOSN5345 88 88 D_lateral AREA=3.125E-016    
M5344 88 430 601 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5343 88 430 446 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5342 446 447 608 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5340 608 601 445 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5339 449 443 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5338 448 430 608 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5337 104 430 601 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5336 608 447 444 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5335 444 601 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M5334 449 443 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D5333 are shorted:
* D5333 88 88 D_lateral AREA=3.125E-016    $ (-1250.5 946.499 -1245.5 946.5)CMOSN5333 88 88 D_lateral AREA=3.125E-016    
M5332 447 460 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5331 88 460 445 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5330 614 460 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M5329 88 503 607 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5328 607 625 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5327 453 449 454 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M5326 88 450 453 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M5325 454 457 458 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M5324 450 451 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5323 447 460 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5322 104 460 448 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5321 104 460 614 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5320 607 503 452 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5319 452 625 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5318 458 449 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M5317 104 450 458 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M5316 104 457 458 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M5315 450 451 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D5314 are shorted:
* D5314 104 104 D_lateral AREA=3.125E-016    $ (-1319 932.499 -1314 932.5)CMOSN5314 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5313 are shorted:
* D5313 88 88 D_lateral AREA=3.125E-016    $ (-1381 946.499 -1376 946.5)CMOSN5313 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5312 are shorted:
* D5312 88 88 D_lateral AREA=3.125E-016    $ (-1335 946 -1334.999 951)CMOSN5312 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5311 are shorted:
* D5311 104 104 D_lateral AREA=3.125E-016    $ (-1328.001 1002.5 -1328 1007.5)CMOSN5311 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5310 are shorted:
* D5310 88 88 D_lateral AREA=3.125E-016    $ (-1329.5 1019.5 -1329.499 1024.5)CMOSN5310 88 88 D_lateral AREA=3.125E-016    
M5309 88 626 617 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M5308 88 460 462 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5307 462 455 618 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5306 455 617 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5305 461 617 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5304 618 614 461 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5303 487 458 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5302 104 626 617 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M5301 456 460 618 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5300 618 455 459 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5299 104 617 456 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5298 455 617 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5297 459 614 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M5296 487 458 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D5295 are shorted:
* D5295 104 104 D_lateral AREA=3.125E-016    $ (-1449.5 932.499 -1444.5 932.5)CMOSN5295 104 104 D_lateral AREA=3.125E-016    
M5294 88 503 626 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5293 626 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5292 626 503 463 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5291 463 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5290 are shorted:
* D5290 88 88 D_lateral AREA=3.125E-016    $ (-1506.5 946 -1506.499 951)CMOSN5290 88 88 D_lateral AREA=3.125E-016    
M5289 88 430 628 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5288 88 430 468 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5287 468 464 629 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5286 464 333 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5285 467 333 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5284 629 628 467 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5283 465 430 629 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5282 104 430 628 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5281 629 464 466 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5280 104 333 465 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5279 464 333 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5278 466 628 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D5277 are shorted:
* D5277 88 88 D_lateral AREA=3.125E-016    $ (-1614 946.499 -1609 946.5)CMOSN5277 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5276 are shorted:
* D5276 104 104 D_lateral AREA=3.125E-016    $ (-1682.5 932.499 -1677.5 932.5)CMOSN5276 104 104 D_lateral AREA=3.125E-016    
M5275 88 469 483 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5274 88 469 475 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5273 475 476 482 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5272 88 333 636 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5271 88 333 474 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5270 474 478 653 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5269 473 652 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5268 653 636 473 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5267 88 503 641 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5266 641 651 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5265 477 469 482 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5264 104 469 483 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5263 482 476 472 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5261 479 333 653 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5260 104 333 636 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5259 653 478 471 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5258 104 652 479 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5257 471 636 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M5256 641 503 470 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5255 470 651 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5254 are shorted:
* D5254 88 88 D_lateral AREA=3.125E-016    $ (-1756.5 1018.499 -1751.5 1018.5)CMOSN5254 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5253 are shorted:
* D5253 88 88 D_lateral AREA=3.125E-016    $ (-1744.5 946.499 -1739.5 946.5)CMOSN5253 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5252 are shorted:
* D5252 88 88 D_lateral AREA=3.125E-016    $ (-1698.5 946 -1698.499 951)CMOSN5252 88 88 D_lateral AREA=3.125E-016    
M5251 476 480 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5250 484 480 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5249 482 483 484 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5248 480 485 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M5246 88 648 652 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M5245 478 652 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5244 88 503 648 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5243 648 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5242 476 480 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5241 104 480 477 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5240 104 483 472 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=187.5f PS=1.25u    
M5239 480 485 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5238 104 648 652 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M5237 478 652 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5236 648 503 481 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5235 104 104 481 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
* Pins of element D5234 are shorted:
* D5234 104 104 D_lateral AREA=3.125E-016    $ (-1825 1004.499 -1820 1004.5)CMOSN5234 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5233 are shorted:
* D5233 88 88 D_lateral AREA=3.125E-016    $ (-1884.5 1018 -1884.499 1023)CMOSN5233 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5232 are shorted:
* D5232 104 104 D_lateral AREA=3.125E-016    $ (-1813 932.499 -1808 932.5)CMOSN5232 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5231 are shorted:
* D5231 88 88 D_lateral AREA=3.125E-016    $ (-1870 946 -1869.999 951)CMOSN5231 88 88 D_lateral AREA=3.125E-016    
M5230 485 487 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5229 485 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5228 485 487 486 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5227 486 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5226 503 489 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M5225 489 657 490 88 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M5224 503 489 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5223 104 657 489 104 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M5222 490 491 88 88 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M5221 506 667 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M5220 88 664 667 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5219 667 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5218 489 491 104 104 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M5217 506 667 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5216 667 664 488 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5215 104 491 488 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
* Pins of element D5214 are shorted:
* D5214 88 88 D_lateral AREA=3.125E-016    $ (-2269.5 946 -2269.499 951)CMOSN5214 88 88 D_lateral AREA=3.125E-016    
M5213 505 498 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5212 88 104 498 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
* Pins of element D5210 are shorted:
* D5210 88 88 D_lateral AREA=3.125E-016    $ (219.5 902 219.501 907)CMOSN5210 88 88 D_lateral AREA=3.125E-016    
M5209 88 493 513 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M5208 493 495 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5207 498 494 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5206 88 494 495 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5205 495 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5204 504 508 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5203 104 493 510 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M5202 493 495 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5201 104 498 505 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5200 497 494 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5199 498 104 497 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5198 495 494 496 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5197 496 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5196 504 508 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D5195 are shorted:
* D5195 88 88 D_lateral AREA=3.125E-016    $ (125.5 857 125.501 862)CMOSN5195 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5194 are shorted:
* D5194 104 104 D_lateral AREA=3.125E-016    $ (126.999 840 127 845)CMOSN5194 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5193 are shorted:
* D5193 88 88 D_lateral AREA=3.125E-016    $ (175 902 175.001 907)CMOSN5193 88 88 D_lateral AREA=3.125E-016    
M5192 543 510 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5191 513 505 514 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M5190 514 516 510 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M5189 88 504 500 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5188 88 504 512 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5187 512 499 710 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5186 499 507 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5185 511 507 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5184 710 500 511 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5183 543 510 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5182 510 505 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M5181 104 516 510 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M5180 501 504 710 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5179 104 504 500 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5178 710 499 509 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5177 104 507 501 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5176 499 507 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5175 509 500 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D5174 are shorted:
* D5174 88 88 D_lateral AREA=3.125E-016    $ (81 902.499 86 902.5)CMOSN5174 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5173 are shorted:
* D5173 104 104 D_lateral AREA=3.125E-016    $ (12.5 888.499 17.5 888.5)CMOSN5173 104 104 D_lateral AREA=3.125E-016    
M5172 516 517 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5171 88 104 517 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5170 517 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5169 516 517 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5168 517 104 519 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5167 519 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5166 are shorted:
* D5166 88 88 D_lateral AREA=3.125E-016    $ (-51.5 902 -51.499 907)CMOSN5166 88 88 D_lateral AREA=3.125E-016    
M5165 523 520 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5164 88 543 520 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5163 520 391 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5162 523 520 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5161 520 543 521 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5160 521 391 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5159 are shorted:
* D5159 88 88 D_lateral AREA=3.125E-016    $ (-144 902 -143.999 907)CMOSN5159 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5158 are shorted:
* D5158 88 88 D_lateral AREA=3.125E-016    $ (-188.5 902 -188.499 907)CMOSN5158 88 88 D_lateral AREA=3.125E-016    
M5157 528 523 529 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M5156 88 524 528 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M5155 529 533 534 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M5154 524 525 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5153 88 391 525 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5152 525 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5151 538 526 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5150 536 538 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M5149 534 523 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M5148 104 524 534 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M5147 104 533 534 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M5146 524 525 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5145 525 391 527 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5144 527 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5143 538 526 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5142 104 538 536 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D5141 are shorted:
* D5141 104 104 D_lateral AREA=3.125E-016    $ (-236.501 840 -236.5 845)CMOSN5141 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5140 are shorted:
* D5140 88 88 D_lateral AREA=3.125E-016    $ (-238 857 -237.999 862)CMOSN5140 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5139 are shorted:
* D5139 88 88 D_lateral AREA=3.125E-016    $ (-282.5 902.499 -277.5 902.5)CMOSN5139 88 88 D_lateral AREA=3.125E-016    
M5138 573 534 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5137 533 541 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5136 88 538 540 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5135 540 530 720 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5134 530 535 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5133 539 535 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5132 720 536 539 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5131 573 534 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5130 533 541 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5129 531 538 720 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5128 720 530 537 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5127 104 535 531 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5126 530 535 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5125 537 536 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D5124 are shorted:
* D5124 104 104 D_lateral AREA=3.125E-016    $ (-351 888.499 -346 888.5)CMOSN5124 104 104 D_lateral AREA=3.125E-016    
M5123 88 543 541 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5122 541 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5121 541 543 545 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5120 545 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5119 are shorted:
* D5119 88 88 D_lateral AREA=3.125E-016    $ (-415 902 -414.999 907)CMOSN5119 88 88 D_lateral AREA=3.125E-016    
M5118 556 548 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5117 555 549 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5116 88 573 549 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5115 549 547 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5114 88 547 548 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5113 548 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5112 556 548 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5111 555 549 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5110 549 573 551 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5109 551 547 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5108 548 547 550 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5107 550 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5106 are shorted:
* D5106 88 88 D_lateral AREA=3.125E-016    $ (-508.5 902 -508.499 907)CMOSN5106 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5105 are shorted:
* D5105 88 88 D_lateral AREA=3.125E-016    $ (-553 902 -552.999 907)CMOSN5105 88 88 D_lateral AREA=3.125E-016    
M5104 599 554 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5103 562 555 563 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M5102 88 556 562 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M5101 563 567 554 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M5100 553 557 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5099 88 553 552 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5098 88 553 561 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5097 561 564 744 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5096 560 569 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5095 744 552 560 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5094 599 554 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5093 554 555 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M5092 104 556 554 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M5091 104 567 554 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M5090 553 557 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5089 565 553 744 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5088 104 553 552 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5087 744 564 559 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5085 559 552 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D5084 are shorted:
* D5084 104 104 D_lateral AREA=3.125E-016    $ (-601.001 840 -601 845)CMOSN5084 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5083 are shorted:
* D5083 88 88 D_lateral AREA=3.125E-016    $ (-602.5 857 -602.499 862)CMOSN5083 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5082 are shorted:
* D5082 88 88 D_lateral AREA=3.125E-016    $ (-647 902.499 -642 902.5)CMOSN5082 88 88 D_lateral AREA=3.125E-016    
M5081 567 570 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5080 88 573 570 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5079 564 569 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5078 567 570 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5076 564 569 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5075 565 569 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
* Pins of element D5074 are shorted:
* D5074 88 88 D_lateral AREA=3.125E-016    $ (-779.5 902 -779.499 907)CMOSN5074 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5073 are shorted:
* D5073 104 104 D_lateral AREA=3.125E-016    $ (-715.5 888.499 -710.5 888.5)CMOSN5073 104 104 D_lateral AREA=3.125E-016    
M5072 570 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5071 588 571 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5070 88 599 571 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5069 571 577 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5068 574 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5067 574 573 570 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5066 588 571 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5065 571 599 572 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5064 572 577 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5063 are shorted:
* D5063 88 88 D_lateral AREA=3.125E-016    $ (-872 902 -871.999 907)CMOSN5063 88 88 D_lateral AREA=3.125E-016    
M5062 581 588 594 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M5061 88 576 581 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M5060 576 578 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5059 88 577 578 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5058 578 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5057 586 579 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5056 587 588 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M5055 104 576 587 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M5054 576 578 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5053 578 577 580 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5052 580 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5051 586 579 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D5050 are shorted:
* D5050 88 88 D_lateral AREA=3.125E-016    $ (-966 857 -965.999 862)CMOSN5050 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5049 are shorted:
* D5049 104 104 D_lateral AREA=3.125E-016    $ (-964.501 840 -964.5 845)CMOSN5049 104 104 D_lateral AREA=3.125E-016    
* Pins of element D5048 are shorted:
* D5048 88 88 D_lateral AREA=3.125E-016    $ (-916.5 902 -916.499 907)CMOSN5048 88 88 D_lateral AREA=3.125E-016    
M5047 625 587 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5046 594 596 587 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M5045 88 586 583 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M5044 88 586 593 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M5043 593 582 770 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M5042 582 590 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5041 592 590 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5040 770 583 592 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M5039 625 587 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5038 104 596 587 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M5037 584 586 770 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M5036 104 586 583 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M5035 770 582 591 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M5034 104 590 584 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5033 582 590 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5032 591 583 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D5031 are shorted:
* D5031 88 88 D_lateral AREA=3.125E-016    $ (-1010.5 902.499 -1005.5 902.5)CMOSN5031 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5030 are shorted:
* D5030 104 104 D_lateral AREA=3.125E-016    $ (-1079 888.499 -1074 888.5)CMOSN5030 104 104 D_lateral AREA=3.125E-016    
M5029 596 597 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5028 88 599 597 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5027 597 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5026 596 597 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5025 597 599 600 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5024 600 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5023 are shorted:
* D5023 88 88 D_lateral AREA=3.125E-016    $ (-1143 902 -1142.999 907)CMOSN5023 88 88 D_lateral AREA=3.125E-016    
M5022 604 602 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5021 88 625 602 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5020 602 608 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5019 88 608 606 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M5018 604 602 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5017 602 625 603 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5016 603 608 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D5015 are shorted:
* D5015 88 88 D_lateral AREA=3.125E-016    $ (-1236 902 -1235.999 907)CMOSN5015 88 88 D_lateral AREA=3.125E-016    
* Pins of element D5014 are shorted:
* D5014 88 88 D_lateral AREA=3.125E-016    $ (-1280.5 902 -1280.499 907)CMOSN5014 88 88 D_lateral AREA=3.125E-016    
M5013 610 604 611 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M5012 88 605 610 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M5011 611 615 616 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M5010 605 606 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5009 606 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M5008 620 607 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M5007 621 620 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M5006 616 604 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M5005 104 605 616 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M5004 104 615 616 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M5003 605 606 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M5002 609 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M5001 606 608 609 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M5000 620 607 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4999 104 620 621 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D4998 are shorted:
* D4998 104 104 D_lateral AREA=3.125E-016    $ (-1328.501 840 -1328.5 845)CMOSN4998 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4997 are shorted:
* D4997 88 88 D_lateral AREA=3.125E-016    $ (-1330 857 -1329.999 862)CMOSN4997 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4996 are shorted:
* D4996 88 88 D_lateral AREA=3.125E-016    $ (-1374.5 902.499 -1369.5 902.5)CMOSN4996 88 88 D_lateral AREA=3.125E-016    
M4995 651 616 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4994 615 624 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4993 88 620 623 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4992 623 612 780 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4991 612 618 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4990 622 618 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4989 780 621 622 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4988 651 616 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4987 615 624 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4986 613 620 780 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4985 780 612 619 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4984 104 618 613 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4983 612 618 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4982 619 621 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D4981 are shorted:
* D4981 104 104 D_lateral AREA=3.125E-016    $ (-1443 888.499 -1438 888.5)CMOSN4981 104 104 D_lateral AREA=3.125E-016    
M4980 88 625 624 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4979 624 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4978 624 625 627 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4977 627 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D4976 are shorted:
* D4976 88 88 D_lateral AREA=3.125E-016    $ (-1507 902 -1506.999 907)CMOSN4976 88 88 D_lateral AREA=3.125E-016    
M4975 640 630 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4974 639 631 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4973 88 651 631 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4972 631 629 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4971 88 629 630 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4970 630 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4969 640 630 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4968 639 631 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4967 631 651 633 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4966 633 629 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4965 630 629 632 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4964 632 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D4963 are shorted:
* D4963 88 88 D_lateral AREA=3.125E-016    $ (-1599.5 902 -1599.499 907)CMOSN4963 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4962 are shorted:
* D4962 88 88 D_lateral AREA=3.125E-016    $ (-1644 902 -1643.999 907)CMOSN4962 88 88 D_lateral AREA=3.125E-016    
M4961 811 638 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4960 645 639 646 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M4959 88 640 645 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M4958 646 649 638 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M4957 637 641 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4956 88 637 634 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M4955 88 637 644 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4954 644 647 805 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4953 643 653 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4952 805 634 643 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4951 811 638 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4950 638 639 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M4949 104 640 638 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M4948 104 649 638 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M4947 637 641 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4946 635 637 805 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4945 104 637 634 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4944 805 647 642 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4943 104 653 635 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4942 642 634 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D4941 are shorted:
* D4941 104 104 D_lateral AREA=3.125E-016    $ (-1692.001 840 -1692 845)CMOSN4941 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4940 are shorted:
* D4940 88 88 D_lateral AREA=3.125E-016    $ (-1693.5 857 -1693.499 862)CMOSN4940 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4939 are shorted:
* D4939 88 88 D_lateral AREA=3.125E-016    $ (-1738 902.499 -1733 902.5)CMOSN4939 88 88 D_lateral AREA=3.125E-016    
M4938 649 650 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4937 88 651 650 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4936 650 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4935 647 653 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4934 649 650 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4933 650 651 654 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4932 654 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4931 647 653 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
* Pins of element D4930 are shorted:
* D4930 88 88 D_lateral AREA=3.125E-016    $ (-1870.5 902 -1870.499 907)CMOSN4930 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4929 are shorted:
* D4929 104 104 D_lateral AREA=3.125E-016    $ (-1806.5 888.499 -1801.5 888.5)CMOSN4929 104 104 D_lateral AREA=3.125E-016    
M4928 88 430 655 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M4927 88 430 662 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4926 662 663 819 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4924 661 668 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4923 819 655 661 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4922 430 658 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M4921 88 482 658 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4920 658 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4919 656 430 819 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4918 104 430 655 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4917 819 663 660 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4916 104 668 656 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4915 660 655 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M4914 430 658 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4913 658 482 659 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4912 659 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D4911 are shorted:
* D4911 88 88 D_lateral AREA=3.125E-016    $ (-2133.5 855.999 -2128.5 856)CMOSN4911 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4910 are shorted:
* D4910 88 88 D_lateral AREA=3.125E-016    $ (-2156.5 900.5 -2156.499 905.5)CMOSN4910 88 88 D_lateral AREA=3.125E-016    
M4909 88 668 663 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4908 668 665 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M4907 88 811 665 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4906 665 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4905 657 666 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M4904 88 664 666 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4903 666 671 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4902 663 668 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4901 668 665 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4900 665 811 670 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4899 670 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4898 657 666 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4897 666 664 669 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4896 669 671 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D4895 are shorted:
* D4895 104 104 D_lateral AREA=3.125E-016    $ (-2202 841.999 -2197 842)CMOSN4895 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4894 are shorted:
* D4894 88 88 D_lateral AREA=3.125E-016    $ (-2261.5 855.5 -2261.499 860.5)CMOSN4894 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4893 are shorted:
* D4893 88 88 D_lateral AREA=3.125E-016    $ (-2240.5 900.5 -2240.499 905.5)CMOSN4893 88 88 D_lateral AREA=3.125E-016    
M4892 671 491 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M4891 671 491 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4890 88 104 822 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
* Pins of element D4888 are shorted:
* D4888 88 88 D_lateral AREA=3.125E-016    $ (219 740.5 219.001 745.5)CMOSN4888 88 88 D_lateral AREA=3.125E-016    
M4887 88 738 673 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M4886 88 738 677 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4885 677 672 824 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4884 672 681 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4883 676 681 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4882 824 673 676 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4881 822 824 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4880 88 824 821 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4879 821 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4878 829 682 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4877 88 683 682 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4876 674 738 824 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4875 104 738 673 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4874 824 672 675 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4873 104 681 674 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4872 672 681 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4871 675 673 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D4868 are shorted:
* D4868 88 88 D_lateral AREA=3.125E-016    $ (204.5 784.999 209.5 785)CMOSN4868 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4867 are shorted:
* D4867 104 104 D_lateral AREA=3.125E-016    $ (136 770.999 141 771)CMOSN4867 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4866 are shorted:
* D4866 88 88 D_lateral AREA=3.125E-016    $ (174.5 740.5 174.501 745.5)CMOSN4866 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4865 are shorted:
* D4865 88 88 D_lateral AREA=3.125E-016    $ (120 784.5 120.001 789.5)CMOSN4865 88 88 D_lateral AREA=3.125E-016    
M4864 88 681 679 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M4863 88 681 689 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4862 689 678 830 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4861 678 691 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4860 688 691 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4859 830 679 688 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4858 682 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4857 88 829 826 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M4856 88 829 687 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4855 687 831 1040 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4854 831 830 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4853 686 830 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4852 1040 826 686 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4851 680 681 830 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4850 104 681 679 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4849 830 678 685 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4848 104 691 680 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4847 678 691 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4846 685 679 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M4845 684 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4844 684 683 682 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D4838 are shorted:
* D4838 88 88 D_lateral AREA=3.125E-016    $ (74 784.999 79 785)CMOSN4838 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4836 are shorted:
* D4836 88 88 D_lateral AREA=3.125E-016    $ (80.5 740.999 85.5 741)CMOSN4836 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4835 are shorted:
* D4835 104 104 D_lateral AREA=3.125E-016    $ (12 726.999 17 727)CMOSN4835 104 104 D_lateral AREA=3.125E-016    
M4834 88 690 691 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M4833 836 838 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4832 88 104 838 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4831 838 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4830 88 683 690 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4829 690 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4828 104 690 691 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M4826 690 683 692 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4825 692 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D4824 are shorted:
* D4824 88 88 D_lateral AREA=3.125E-016    $ (-52 740.5 -51.999 745.5)CMOSN4824 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4823 are shorted:
* D4823 104 104 D_lateral AREA=3.125E-016    $ (5.5 770.999 10.5 771)CMOSN4823 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4822 are shorted:
* D4822 88 88 D_lateral AREA=3.125E-016    $ (-51.5 784.5 -51.499 789.5)CMOSN4822 88 88 D_lateral AREA=3.125E-016    
M4821 88 738 699 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M4820 88 738 693 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4819 693 696 698 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4818 88 856 839 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4817 839 698 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4816 694 738 698 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4815 104 738 699 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D4813 are shorted:
* D4813 88 88 D_lateral AREA=3.125E-016    $ (-159 784.999 -154 785)CMOSN4813 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4812 are shorted:
* D4812 88 88 D_lateral AREA=3.125E-016    $ (-144.5 740.5 -144.499 745.5)CMOSN4812 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4811 are shorted:
* D4811 88 88 D_lateral AREA=3.125E-016    $ (-189 740.5 -188.999 745.5)CMOSN4811 88 88 D_lateral AREA=3.125E-016    
M4810 696 710 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4809 700 710 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4808 698 699 700 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4807 88 698 843 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4806 843 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4805 851 844 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4803 88 683 844 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4802 844 856 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4801 704 851 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M4800 697 696 698 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=1.84375p PS=4.375u    
M4799 696 710 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4798 104 710 694 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4797 697 699 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M4795 104 710 702 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4794 844 683 695 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4793 695 856 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D4791 are shorted:
* D4791 104 104 D_lateral AREA=3.125E-016    $ (-227.5 770.999 -222.5 771)CMOSN4791 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4790 are shorted:
* D4790 88 88 D_lateral AREA=3.125E-016    $ (-289.5 784.999 -284.5 785)CMOSN4790 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4789 are shorted:
* D4789 88 88 D_lateral AREA=3.125E-016    $ (-243.5 784.5 -243.499 789.5)CMOSN4789 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4788 are shorted:
* D4788 88 88 D_lateral AREA=3.125E-016    $ (-283 740.999 -278 741)CMOSN4788 88 88 D_lateral AREA=3.125E-016    
M4787 88 711 712 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M4786 849 855 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4785 702 710 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M4784 88 710 709 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4783 709 701 852 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4782 701 712 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4781 708 712 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4780 852 702 708 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4779 88 851 707 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4778 707 853 1059 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4777 853 852 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4776 706 852 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4775 1059 704 706 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4774 104 711 712 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M4772 703 710 852 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4771 852 701 705 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4770 104 712 703 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4769 701 712 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4768 705 702 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D4763 are shorted:
* D4763 104 104 D_lateral AREA=3.125E-016    $ (-358 770.999 -353 771)CMOSN4763 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4762 are shorted:
* D4762 104 104 D_lateral AREA=3.125E-016    $ (-351.5 726.999 -346.5 727)CMOSN4762 104 104 D_lateral AREA=3.125E-016    
M4761 88 856 855 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4760 855 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4759 88 683 711 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4758 711 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4757 711 683 713 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4756 713 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D4755 are shorted:
* D4755 88 88 D_lateral AREA=3.125E-016    $ (-415.5 740.5 -415.499 745.5)CMOSN4755 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4754 are shorted:
* D4754 88 88 D_lateral AREA=3.125E-016    $ (-415 784.5 -414.999 789.5)CMOSN4754 88 88 D_lateral AREA=3.125E-016    
M4753 88 738 715 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M4752 88 738 719 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4751 719 714 861 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4750 714 720 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4749 718 720 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4748 861 715 718 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4747 88 879 859 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4746 859 861 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4745 88 861 858 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4744 858 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4743 716 738 861 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4742 104 738 715 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4741 861 714 717 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4740 104 720 716 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4739 714 720 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4738 717 715 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D4737 are shorted:
* D4737 88 88 D_lateral AREA=3.125E-016    $ (-523.5 784.999 -518.5 785)CMOSN4737 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4735 are shorted:
* D4735 88 88 D_lateral AREA=3.125E-016    $ (-509 740.5 -508.999 745.5)CMOSN4735 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4734 are shorted:
* D4734 88 88 D_lateral AREA=3.125E-016    $ (-553.5 740.5 -553.499 745.5)CMOSN4734 88 88 D_lateral AREA=3.125E-016    
M4733 867 869 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4732 88 720 729 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M4731 88 720 725 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4730 725 726 875 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4728 88 683 869 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4727 869 879 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4726 88 867 863 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M4725 88 867 724 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4724 724 872 1102 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4723 723 875 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4722 1102 863 723 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4720 727 720 875 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4719 104 720 729 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4718 875 726 722 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4717 722 729 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M4716 869 683 721 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4715 721 879 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D4709 are shorted:
* D4709 104 104 D_lateral AREA=3.125E-016    $ (-592 770.999 -587 771)CMOSN4709 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4708 are shorted:
* D4708 88 88 D_lateral AREA=3.125E-016    $ (-654 784.999 -649 785)CMOSN4708 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4707 are shorted:
* D4707 88 88 D_lateral AREA=3.125E-016    $ (-608 784.5 -607.999 789.5)CMOSN4707 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4706 are shorted:
* D4706 88 88 D_lateral AREA=3.125E-016    $ (-647.5 740.999 -642.5 741)CMOSN4706 88 88 D_lateral AREA=3.125E-016    
M4705 88 731 728 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M4704 874 876 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4703 88 879 876 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4702 726 728 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4701 730 728 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4700 730 729 875 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4699 88 683 731 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4698 872 875 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4697 104 731 728 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M4695 726 728 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4694 104 728 727 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D4691 are shorted:
* D4691 88 88 D_lateral AREA=3.125E-016    $ (-780 740.5 -779.999 745.5)CMOSN4691 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4690 are shorted:
* D4690 104 104 D_lateral AREA=3.125E-016    $ (-722.5 770.999 -717.5 771)CMOSN4690 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4689 are shorted:
* D4689 88 88 D_lateral AREA=3.125E-016    $ (-779.5 784.5 -779.499 789.5)CMOSN4689 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4688 are shorted:
* D4688 104 104 D_lateral AREA=3.125E-016    $ (-716 726.999 -711 727)CMOSN4688 104 104 D_lateral AREA=3.125E-016    
M4687 876 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4686 731 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4685 734 738 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M4684 88 897 877 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4682 732 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4681 732 683 731 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4680 104 738 734 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D4679 are shorted:
* D4679 88 88 D_lateral AREA=3.125E-016    $ (-887 784.999 -882 785)CMOSN4679 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4678 are shorted:
* D4678 88 88 D_lateral AREA=3.125E-016    $ (-872.5 740.5 -872.499 745.5)CMOSN4678 88 88 D_lateral AREA=3.125E-016    
M4677 88 738 740 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4676 740 733 885 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4675 733 744 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4674 739 744 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4673 885 734 739 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4672 88 885 877 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4671 88 885 882 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4670 882 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4669 890 883 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4668 88 683 883 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4667 883 897 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4666 735 738 885 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4665 885 733 737 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4664 104 744 735 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4663 733 744 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4662 737 734 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M4660 883 683 736 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4659 736 897 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D4658 are shorted:
* D4658 104 104 D_lateral AREA=3.125E-016    $ (-955.5 770.999 -950.5 771)CMOSN4658 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4657 are shorted:
* D4657 88 88 D_lateral AREA=3.125E-016    $ (-917 740.5 -916.999 745.5)CMOSN4657 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4656 are shorted:
* D4656 88 88 D_lateral AREA=3.125E-016    $ (-971.5 784.5 -971.499 789.5)CMOSN4656 88 88 D_lateral AREA=3.125E-016    
M4655 88 744 742 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M4654 88 744 749 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4653 749 741 891 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4652 741 751 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4651 748 751 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4650 891 742 748 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4649 88 890 887 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M4648 88 890 747 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4647 747 892 1146 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4646 892 891 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4645 746 891 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4644 1146 887 746 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4643 743 744 891 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4642 104 744 742 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4641 891 741 745 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4640 104 751 743 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4639 741 751 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4638 745 742 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D4632 are shorted:
* D4632 88 88 D_lateral AREA=3.125E-016    $ (-1017.5 784.999 -1012.5 785)CMOSN4632 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4631 are shorted:
* D4631 104 104 D_lateral AREA=3.125E-016    $ (-1086 770.999 -1081 771)CMOSN4631 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4630 are shorted:
* D4630 88 88 D_lateral AREA=3.125E-016    $ (-1011 740.999 -1006 741)CMOSN4630 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4629 are shorted:
* D4629 104 104 D_lateral AREA=3.125E-016    $ (-1079.5 726.999 -1074.5 727)CMOSN4629 104 104 D_lateral AREA=3.125E-016    
M4628 88 750 751 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M4627 896 899 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4626 88 897 899 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4625 899 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4624 88 683 750 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4623 750 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4622 104 750 751 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M4620 750 683 752 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4619 752 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D4618 are shorted:
* D4618 88 88 D_lateral AREA=3.125E-016    $ (-1143.5 740.5 -1143.499 745.5)CMOSN4618 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4617 are shorted:
* D4617 88 88 D_lateral AREA=3.125E-016    $ (-1143 784.5 -1142.999 789.5)CMOSN4617 88 88 D_lateral AREA=3.125E-016    
M4616 88 738 759 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M4615 88 738 753 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4614 753 754 758 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4613 88 917 900 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4612 900 758 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4611 755 738 758 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4610 104 738 759 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4609 758 754 757 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
* Pins of element D4608 are shorted:
* D4608 88 88 D_lateral AREA=3.125E-016    $ (-1258.5 784.999 -1253.5 785)CMOSN4608 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4607 are shorted:
* D4607 88 88 D_lateral AREA=3.125E-016    $ (-1244 740.5 -1243.999 745.5)CMOSN4607 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4606 are shorted:
* D4606 88 88 D_lateral AREA=3.125E-016    $ (-1288.5 740.5 -1288.499 745.5)CMOSN4606 88 88 D_lateral AREA=3.125E-016    
M4605 754 770 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4604 760 770 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4603 758 759 760 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4602 88 758 904 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4601 904 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4600 912 905 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4598 88 683 905 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4597 905 917 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4596 764 912 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M4595 754 770 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4594 104 770 755 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4593 757 759 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M4591 104 770 762 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4590 905 683 756 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4589 756 917 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D4587 are shorted:
* D4587 104 104 D_lateral AREA=3.125E-016    $ (-1327 770.999 -1322 771)CMOSN4587 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4586 are shorted:
* D4586 88 88 D_lateral AREA=3.125E-016    $ (-1389 784.999 -1384 785)CMOSN4586 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4585 are shorted:
* D4585 88 88 D_lateral AREA=3.125E-016    $ (-1343 784.5 -1342.999 789.5)CMOSN4585 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4584 are shorted:
* D4584 88 88 D_lateral AREA=3.125E-016    $ (-1382.5 740.999 -1377.5 741)CMOSN4584 88 88 D_lateral AREA=3.125E-016    
M4583 88 771 772 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M4582 910 916 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4581 762 770 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M4580 88 770 769 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4579 769 761 913 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4578 761 772 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4577 768 772 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4576 913 762 768 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4575 88 912 767 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4574 767 914 1165 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4573 914 913 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4572 766 913 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4571 1165 764 766 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4570 104 771 772 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M4568 763 770 913 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4567 913 761 765 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4566 104 772 763 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4565 761 772 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4564 765 762 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D4559 are shorted:
* D4559 104 104 D_lateral AREA=3.125E-016    $ (-1457.5 770.999 -1452.5 771)CMOSN4559 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4558 are shorted:
* D4558 104 104 D_lateral AREA=3.125E-016    $ (-1451 726.999 -1446 727)CMOSN4558 104 104 D_lateral AREA=3.125E-016    
M4557 88 917 916 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4556 916 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4555 88 683 771 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4554 771 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4553 771 683 773 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4552 773 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D4551 are shorted:
* D4551 88 88 D_lateral AREA=3.125E-016    $ (-1515 740.5 -1514.999 745.5)CMOSN4551 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4550 are shorted:
* D4550 88 88 D_lateral AREA=3.125E-016    $ (-1514.5 784.5 -1514.499 789.5)CMOSN4550 88 88 D_lateral AREA=3.125E-016    
M4549 88 738 775 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M4548 88 738 779 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4547 779 774 922 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4546 774 780 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4545 778 780 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4544 922 775 778 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4543 88 937 920 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4542 920 922 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4541 88 922 919 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4540 919 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4539 776 738 922 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4538 104 738 775 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4537 922 774 777 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4536 104 780 776 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4535 774 780 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4534 777 775 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D4533 are shorted:
* D4533 88 88 D_lateral AREA=3.125E-016    $ (-1627 784.999 -1622 785)CMOSN4533 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4531 are shorted:
* D4531 88 88 D_lateral AREA=3.125E-016    $ (-1612.5 740.5 -1612.499 745.5)CMOSN4531 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4530 are shorted:
* D4530 88 88 D_lateral AREA=3.125E-016    $ (-1657 740.5 -1656.999 745.5)CMOSN4530 88 88 D_lateral AREA=3.125E-016    
M4529 927 929 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4528 88 780 790 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M4527 88 780 784 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4526 784 785 789 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4525 88 683 929 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4524 929 937 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4523 88 927 924 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M4522 88 927 783 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4521 783 932 1206 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4519 1206 924 782 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4517 786 780 789 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4516 104 780 790 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4515 789 785 788 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4514 929 683 781 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4513 781 937 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D4508 are shorted:
* D4508 104 104 D_lateral AREA=3.125E-016    $ (-1695.5 770.999 -1690.5 771)CMOSN4508 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4507 are shorted:
* D4507 88 88 D_lateral AREA=3.125E-016    $ (-1757.5 784.999 -1752.5 785)CMOSN4507 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4506 are shorted:
* D4506 88 88 D_lateral AREA=3.125E-016    $ (-1711.5 784.5 -1711.499 789.5)CMOSN4506 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4505 are shorted:
* D4505 88 88 D_lateral AREA=3.125E-016    $ (-1751 740.999 -1746 741)CMOSN4505 88 88 D_lateral AREA=3.125E-016    
M4504 88 792 787 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M4503 934 936 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4501 785 787 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4500 791 787 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4499 789 790 791 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4497 932 789 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4496 88 789 782 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4495 104 792 787 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M4493 785 787 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4492 104 787 786 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4491 788 790 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D4489 are shorted:
* D4489 88 88 D_lateral AREA=3.125E-016    $ (-1883.5 740.5 -1883.499 745.5)CMOSN4489 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4488 are shorted:
* D4488 104 104 D_lateral AREA=3.125E-016    $ (-1826 770.999 -1821 771)CMOSN4488 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4487 are shorted:
* D4487 88 88 D_lateral AREA=3.125E-016    $ (-1883 784.5 -1882.999 789.5)CMOSN4487 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4486 are shorted:
* D4486 104 104 D_lateral AREA=3.125E-016    $ (-1819.5 726.999 -1814.5 727)CMOSN4486 104 104 D_lateral AREA=3.125E-016    
M4485 88 956 799 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4484 936 937 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4483 936 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4482 792 683 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4481 792 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4480 104 738 795 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4479 792 683 793 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4478 793 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D4477 are shorted:
* D4477 88 88 D_lateral AREA=3.125E-016    $ (-1990.5 784.999 -1985.5 785)CMOSN4477 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4476 are shorted:
* D4476 88 88 D_lateral AREA=3.125E-016    $ (-1976 740.5 -1975.999 745.5)CMOSN4476 88 88 D_lateral AREA=3.125E-016    
M4475 88 738 795 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M4474 88 738 801 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4473 801 794 944 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4472 794 805 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4471 800 805 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4470 944 795 800 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4469 799 944 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4468 88 944 940 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4467 940 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4466 950 941 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4465 88 683 941 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4463 796 738 944 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4462 944 794 798 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4461 104 805 796 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4460 794 805 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4459 798 795 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M4457 941 683 797 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
* Pins of element D4455 are shorted:
* D4455 104 104 D_lateral AREA=3.125E-016    $ (-2059 770.999 -2054 771)CMOSN4455 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4454 are shorted:
* D4454 88 88 D_lateral AREA=3.125E-016    $ (-2020.5 740.5 -2020.499 745.5)CMOSN4454 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4453 are shorted:
* D4453 88 88 D_lateral AREA=3.125E-016    $ (-2075 784.5 -2074.999 789.5)CMOSN4453 88 88 D_lateral AREA=3.125E-016    
M4452 88 805 803 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M4451 88 805 810 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4450 810 802 951 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4449 802 813 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4448 809 813 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4447 951 803 809 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4446 88 956 941 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4445 88 950 946 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M4444 88 950 808 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4443 808 952 1241 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4442 952 951 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4441 807 951 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4440 1241 946 807 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4439 804 805 951 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4438 104 805 803 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4437 951 802 806 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4436 104 813 804 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4435 802 813 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4434 806 803 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M4433 104 956 797 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
* Pins of element D4427 are shorted:
* D4427 88 88 D_lateral AREA=3.125E-016    $ (-2121 784.999 -2116 785)CMOSN4427 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4426 are shorted:
* D4426 104 104 D_lateral AREA=3.125E-016    $ (-2189.5 770.999 -2184.5 771)CMOSN4426 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4425 are shorted:
* D4425 88 88 D_lateral AREA=3.125E-016    $ (-2114.5 740.999 -2109.5 741)CMOSN4425 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4424 are shorted:
* D4424 104 104 D_lateral AREA=3.125E-016    $ (-2183 726.999 -2178 727)CMOSN4424 104 104 D_lateral AREA=3.125E-016    
M4423 88 812 813 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M4422 955 958 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4421 88 956 958 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4420 958 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4419 88 683 812 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4418 812 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4417 104 812 813 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M4415 812 683 814 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4414 814 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D4413 are shorted:
* D4413 88 88 D_lateral AREA=3.125E-016    $ (-2247 740.5 -2246.999 745.5)CMOSN4413 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4412 are shorted:
* D4412 88 88 D_lateral AREA=3.125E-016    $ (-2246.5 784.5 -2246.499 789.5)CMOSN4412 88 88 D_lateral AREA=3.125E-016    
M4411 738 964 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M4410 88 819 964 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4409 964 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4408 683 815 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M4407 816 491 88 88 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M4406 815 962 816 88 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M4405 962 971 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M4404 683 815 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4403 815 491 104 104 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M4402 104 962 815 104 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
* Pins of element D4401 are shorted:
* D4401 88 88 D_lateral AREA=3.125E-016    $ (-2527.5 739 -2527.499 744)CMOSN4401 88 88 D_lateral AREA=3.125E-016    
M4400 88 973 971 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4399 971 972 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4398 972 491 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M4397 681 817 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M4396 88 973 817 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4395 817 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4394 681 817 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4393 817 973 818 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4392 818 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D4391 are shorted:
* D4391 88 88 D_lateral AREA=3.125E-016    $ (-2611.5 739 -2611.499 744)CMOSN4391 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4390 are shorted:
* D4390 88 88 D_lateral AREA=3.125E-016    $ (-2640.5 784.5 -2640.499 789.5)CMOSN4390 88 88 D_lateral AREA=3.125E-016    
M4380 88 820 834 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M4379 820 821 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4378 88 822 828 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4377 104 820 833 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M4376 820 821 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4375 104 822 828 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4374 822 104 825 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4373 825 824 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4372 821 824 823 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4371 823 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4370 829 682 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D4368 are shorted:
* D4368 88 88 D_lateral AREA=3.125E-016    $ (125 695.5 125.001 700.5)CMOSN4368 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4367 are shorted:
* D4367 104 104 D_lateral AREA=3.125E-016    $ (126.499 678.5 126.5 683.5)CMOSN4367 104 104 D_lateral AREA=3.125E-016    
M4359 856 833 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4358 834 828 835 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M4357 835 836 833 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M4356 856 833 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4355 833 828 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M4354 104 836 833 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M4353 1040 831 832 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4352 831 830 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4351 832 826 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M4350 104 830 827 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4349 827 829 1040 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4348 104 829 826 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4344 836 838 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4343 838 104 837 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4342 837 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4337 841 839 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4336 841 839 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4335 839 856 840 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4334 840 698 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4327 846 841 847 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M4326 88 842 846 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M4325 847 849 850 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M4324 842 843 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4323 850 841 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M4322 104 842 850 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M4321 104 849 850 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M4320 842 843 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4319 843 698 845 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4318 845 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4317 851 844 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4316 104 851 704 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D4314 are shorted:
* D4314 104 104 D_lateral AREA=3.125E-016    $ (-237.001 678.5 -237 683.5)CMOSN4314 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4313 are shorted:
* D4313 88 88 D_lateral AREA=3.125E-016    $ (-238.5 695.5 -238.499 700.5)CMOSN4313 88 88 D_lateral AREA=3.125E-016    
M4305 879 850 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4304 879 850 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4303 849 855 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4302 1059 853 854 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4301 853 852 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4300 854 704 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M4299 104 852 848 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4298 848 851 1059 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4295 855 856 857 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4294 857 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4286 866 858 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4285 865 859 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4284 866 858 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4283 865 859 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4282 859 879 862 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4281 862 861 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4280 858 861 860 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4279 860 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4272 897 864 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4271 870 865 871 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M4270 88 866 870 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M4269 871 874 864 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M4268 897 864 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4267 864 865 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M4266 104 866 864 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M4265 104 874 864 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M4264 867 869 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4263 1102 872 868 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4262 868 863 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M4260 873 867 1102 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4259 104 867 863 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D4257 are shorted:
* D4257 104 104 D_lateral AREA=3.125E-016    $ (-601.501 678.5 -601.5 683.5)CMOSN4257 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4256 are shorted:
* D4256 88 88 D_lateral AREA=3.125E-016    $ (-603 695.5 -602.999 700.5)CMOSN4256 88 88 D_lateral AREA=3.125E-016    
M4250 874 876 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4248 872 875 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4247 873 875 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4243 894 877 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4242 880 879 876 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4241 880 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4240 894 877 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4239 877 897 878 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4230 886 894 895 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M4229 88 881 886 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M4228 881 882 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4226 104 881 889 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M4225 881 882 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4224 104 885 878 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4223 882 885 884 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4222 884 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4221 890 883 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D4219 are shorted:
* D4219 88 88 D_lateral AREA=3.125E-016    $ (-966.5 695.5 -966.499 700.5)CMOSN4219 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4218 are shorted:
* D4218 104 104 D_lateral AREA=3.125E-016    $ (-965.001 678.5 -965 683.5)CMOSN4218 104 104 D_lateral AREA=3.125E-016    
M4211 917 889 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4210 895 896 889 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M4209 917 889 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4208 104 896 889 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M4207 104 894 889 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=1.15625p PS=3.5u    
M4206 1146 892 893 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4205 892 891 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4204 893 887 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M4203 104 891 888 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4202 888 890 1146 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4201 104 890 887 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4197 896 899 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4196 899 897 898 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4195 898 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4190 902 900 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4189 902 900 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4188 900 917 901 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4187 901 758 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4180 907 902 908 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M4179 88 903 907 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M4178 908 910 911 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M4177 903 904 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4176 911 902 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M4175 104 903 911 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M4174 104 910 911 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M4173 903 904 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4172 904 758 906 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4171 906 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4170 912 905 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4169 104 912 764 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D4167 are shorted:
* D4167 104 104 D_lateral AREA=3.125E-016    $ (-1336.501 678.5 -1336.5 683.5)CMOSN4167 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4166 are shorted:
* D4166 88 88 D_lateral AREA=3.125E-016    $ (-1338 695.5 -1337.999 700.5)CMOSN4166 88 88 D_lateral AREA=3.125E-016    
M4158 937 911 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4157 937 911 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4156 910 916 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4155 1165 914 915 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4154 914 913 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4153 915 764 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M4152 104 913 909 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4151 909 912 1165 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4148 916 917 918 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4147 918 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4139 926 919 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4138 925 920 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4137 926 919 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4136 925 920 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4135 920 937 923 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4134 923 922 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4133 919 922 921 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4132 921 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4126 956 935 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4125 930 925 931 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M4124 88 926 930 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M4123 931 934 935 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M4122 956 935 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4121 935 925 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M4120 104 926 935 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M4119 104 934 935 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M4118 927 929 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4117 1206 932 928 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4116 928 924 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M4115 933 927 1206 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4114 104 927 924 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D4112 are shorted:
* D4112 104 104 D_lateral AREA=3.125E-016    $ (-1705.001 678.5 -1705 683.5)CMOSN4112 104 104 D_lateral AREA=3.125E-016    
* Pins of element D4111 are shorted:
* D4111 88 88 D_lateral AREA=3.125E-016    $ (-1706.5 695.5 -1706.499 700.5)CMOSN4111 88 88 D_lateral AREA=3.125E-016    
M4105 934 936 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4104 932 789 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4103 104 789 933 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4099 949 799 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4098 949 799 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4097 799 956 943 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4096 936 937 938 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4095 938 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4086 88 939 945 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M4085 939 940 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4083 104 939 948 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M4082 939 940 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4081 943 944 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4080 940 944 942 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4079 942 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4078 950 941 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D4076 are shorted:
* D4076 88 88 D_lateral AREA=3.125E-016    $ (-2070 695.5 -2069.999 700.5)CMOSN4076 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4075 are shorted:
* D4075 104 104 D_lateral AREA=3.125E-016    $ (-2068.501 678.5 -2068.5 683.5)CMOSN4075 104 104 D_lateral AREA=3.125E-016    
M4067 969 948 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M4066 954 949 945 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.125p PS=3.75u    
M4065 954 955 948 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M4064 969 948 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4063 104 949 948 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=1.15625p PS=3.5u    
M4062 104 955 948 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M4061 1241 952 953 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4060 952 951 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4059 953 946 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M4058 104 951 947 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4057 947 950 1241 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4056 104 950 946 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4052 955 958 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M4051 958 956 957 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4050 957 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4039 88 738 960 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M4038 88 738 967 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M4037 967 959 976 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M4036 959 968 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4035 966 968 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4034 976 960 966 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M4026 961 738 976 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M4025 104 738 960 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4024 976 959 965 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M4023 104 968 961 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4022 959 968 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M4021 965 960 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M4020 738 964 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4019 964 819 963 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4018 963 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4017 962 971 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D4016 are shorted:
* D4016 88 88 D_lateral AREA=3.125E-016    $ (-2504.5 694.499 -2499.5 694.5)CMOSN4016 88 88 D_lateral AREA=3.125E-016    
* Pins of element D4015 are shorted:
* D4015 104 104 D_lateral AREA=3.125E-016    $ (-2573 680.499 -2568 680.5)CMOSN4015 104 104 D_lateral AREA=3.125E-016    
M4014 968 970 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M4013 88 969 970 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M4012 970 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M4009 968 970 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M4008 970 969 975 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4007 975 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4006 971 973 974 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M4005 974 972 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M4004 972 491 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D4003 are shorted:
* D4003 88 88 D_lateral AREA=3.125E-016    $ (-2632.5 694 -2632.499 699)CMOSN4003 88 88 D_lateral AREA=3.125E-016    
M3993 88 104 1276 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
* Pins of element D3991 are shorted:
* D3991 88 88 D_lateral AREA=3.125E-016    $ (218.5 578 218.501 583)CMOSN3991 88 88 D_lateral AREA=3.125E-016    
M3990 88 1093 978 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3989 88 1093 985 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3988 985 977 980 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3987 977 994 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3986 88 994 984 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3985 980 978 984 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3984 88 1277 1004 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M3983 1277 1275 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3982 88 1276 1286 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3981 1276 980 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3980 88 980 1275 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3979 1275 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3978 992 993 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3977 88 997 993 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3976 979 1093 980 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3975 104 1093 978 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3974 980 977 983 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3973 104 994 979 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3972 977 994 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3971 983 978 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3970 982 980 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3969 1276 104 982 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3968 1275 980 981 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3967 981 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3966 992 993 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D3965 are shorted:
* D3965 88 88 D_lateral AREA=3.125E-016    $ (204 622.499 209 622.5)CMOSN3965 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3964 are shorted:
* D3964 104 104 D_lateral AREA=3.125E-016    $ (135.5 608.499 140.5 608.5)CMOSN3964 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3963 are shorted:
* D3963 88 88 D_lateral AREA=3.125E-016    $ (124.5 533 124.501 538)CMOSN3963 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3962 are shorted:
* D3962 88 88 D_lateral AREA=3.125E-016    $ (174 578 174.001 583)CMOSN3962 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3961 are shorted:
* D3961 88 88 D_lateral AREA=3.125E-016    $ (119.5 622 119.501 627)CMOSN3961 88 88 D_lateral AREA=3.125E-016    
M3960 1042 1285 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3959 1004 1286 1005 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M3958 1005 1007 1285 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M3957 88 994 987 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3956 88 994 1003 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3955 1003 986 995 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3954 986 1006 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3953 88 1006 1002 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3952 995 987 1002 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3951 993 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3950 88 992 990 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3949 88 992 1001 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3948 1001 989 1295 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3947 989 995 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3946 1000 995 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3945 1295 990 1000 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3944 988 994 995 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3943 104 994 987 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3942 995 986 999 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3941 104 1006 988 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3940 986 1006 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3939 999 987 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3938 998 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3937 993 997 998 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3936 991 992 1295 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3935 104 992 990 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3934 1295 989 996 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3933 104 995 991 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3932 989 995 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3931 996 990 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D3930 are shorted:
* D3930 88 88 D_lateral AREA=3.125E-016    $ (73.5 622.499 78.5 622.5)CMOSN3930 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3928 are shorted:
* D3928 88 88 D_lateral AREA=3.125E-016    $ (80 578.499 85 578.5)CMOSN3928 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3927 are shorted:
* D3927 104 104 D_lateral AREA=3.125E-016    $ (11.5 564.499 16.5 564.5)CMOSN3927 104 104 D_lateral AREA=3.125E-016    
M3926 88 1009 1006 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M3925 1007 1008 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3924 88 104 1008 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3923 1008 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3922 88 997 1009 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3921 1009 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3920 104 1009 1006 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M3919 1007 1008 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3918 1008 104 1011 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3917 1011 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3916 1009 997 1010 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3915 1010 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D3914 are shorted:
* D3914 88 88 D_lateral AREA=3.125E-016    $ (-52.5 578 -52.499 583)CMOSN3914 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3913 are shorted:
* D3913 104 104 D_lateral AREA=3.125E-016    $ (5 608.499 10 608.5)CMOSN3913 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3912 are shorted:
* D3912 88 88 D_lateral AREA=3.125E-016    $ (-52 622 -51.999 627)CMOSN3912 88 88 D_lateral AREA=3.125E-016    
M3911 88 1093 1023 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3910 88 1093 1013 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3909 1013 1018 1022 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3908 1299 1296 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3907 88 1042 1296 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3906 1296 1022 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3905 1014 1093 1022 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3904 104 1093 1023 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3902 1296 1042 1012 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3901 1012 1022 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D3900 are shorted:
* D3900 88 88 D_lateral AREA=3.125E-016    $ (-159.5 622.499 -154.5 622.5)CMOSN3900 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3899 are shorted:
* D3899 88 88 D_lateral AREA=3.125E-016    $ (-145 578 -144.999 583)CMOSN3899 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3898 are shorted:
* D3898 88 88 D_lateral AREA=3.125E-016    $ (-189.5 578 -189.499 583)CMOSN3898 88 88 D_lateral AREA=3.125E-016    
M3897 1018 1040 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3896 88 1040 1024 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3895 1022 1023 1024 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3894 1020 1299 1021 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M3893 88 1301 1020 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M3892 1021 1031 1311 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M3891 1301 1300 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3890 88 1022 1300 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3889 1300 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3888 1034 1015 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3886 88 997 1015 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3885 1015 1042 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3884 1029 1034 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M3883 1019 1018 1022 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=1.84375p PS=4.375u    
M3882 1018 1040 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3881 104 1040 1014 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3880 1019 1023 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3879 1300 1022 1017 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3878 1017 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3877 1034 1015 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3876 104 1040 1026 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3875 1015 997 1016 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3874 1016 1042 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3873 104 1034 1029 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D3872 are shorted:
* D3872 104 104 D_lateral AREA=3.125E-016    $ (-228 608.499 -223 608.5)CMOSN3872 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3871 are shorted:
* D3871 88 88 D_lateral AREA=3.125E-016    $ (-239 533 -238.999 538)CMOSN3871 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3870 are shorted:
* D3870 88 88 D_lateral AREA=3.125E-016    $ (-290 622.499 -285 622.5)CMOSN3870 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3869 are shorted:
* D3869 88 88 D_lateral AREA=3.125E-016    $ (-244 622 -243.999 627)CMOSN3869 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3868 are shorted:
* D3868 88 88 D_lateral AREA=3.125E-016    $ (-283.5 578.499 -278.5 578.5)CMOSN3868 88 88 D_lateral AREA=3.125E-016    
M3867 88 1044 1041 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M3866 1081 1311 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3865 1031 1043 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3864 1026 1040 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M3863 88 1040 1039 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3862 1039 1025 1032 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3861 1025 1041 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3860 88 1041 1038 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3859 1032 1026 1038 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3858 88 1034 1037 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3857 1037 1028 1317 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3856 1028 1032 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3855 1036 1032 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3854 1317 1029 1036 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3853 104 1044 1041 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M3852 1031 1043 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3851 1027 1040 1032 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3850 1032 1025 1035 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3849 104 1041 1027 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3848 1025 1041 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3847 1035 1026 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3846 1030 1034 1317 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3845 1317 1028 1033 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3844 104 1032 1030 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3843 1028 1032 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3842 1033 1029 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D3841 are shorted:
* D3841 104 104 D_lateral AREA=3.125E-016    $ (-358.5 608.499 -353.5 608.5)CMOSN3841 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3840 are shorted:
* D3840 104 104 D_lateral AREA=3.125E-016    $ (-352 564.499 -347 564.5)CMOSN3840 104 104 D_lateral AREA=3.125E-016    
M3839 88 1042 1043 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3838 1043 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3837 88 997 1044 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3836 1044 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3835 1043 1042 1046 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3834 1046 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3833 1044 997 1045 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3832 1045 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D3831 are shorted:
* D3831 88 88 D_lateral AREA=3.125E-016    $ (-416 578 -415.999 583)CMOSN3831 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3830 are shorted:
* D3830 88 88 D_lateral AREA=3.125E-016    $ (-415.5 622 -415.499 627)CMOSN3830 88 88 D_lateral AREA=3.125E-016    
M3829 88 1093 1048 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3828 88 1093 1055 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3827 1055 1047 1050 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3826 1047 1059 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3825 88 1059 1054 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3824 1050 1048 1054 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3823 1329 1322 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3822 1328 1323 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3821 88 1081 1323 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3820 1323 1050 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3819 88 1050 1322 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3818 1322 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3817 1049 1093 1050 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3816 104 1093 1048 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3815 1050 1047 1053 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3814 104 1059 1049 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3813 1047 1059 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3812 1053 1048 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3811 1323 1081 1052 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3810 1052 1050 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3809 1322 1050 1051 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3808 1051 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D3807 are shorted:
* D3807 88 88 D_lateral AREA=3.125E-016    $ (-524 622.499 -519 622.5)CMOSN3807 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3805 are shorted:
* D3805 88 88 D_lateral AREA=3.125E-016    $ (-509.5 578 -509.499 583)CMOSN3805 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3804 are shorted:
* D3804 88 88 D_lateral AREA=3.125E-016    $ (-554 578 -553.999 583)CMOSN3804 88 88 D_lateral AREA=3.125E-016    
M3803 1112 1327 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3802 1066 1328 1067 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M3801 88 1329 1066 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M3800 1067 1073 1327 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M3799 1057 1058 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3798 88 1059 1075 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3797 88 1059 1065 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3796 1065 1068 1074 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3794 88 997 1058 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3793 1058 1081 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3792 88 1057 1056 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3791 88 1057 1064 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3790 1064 1070 1339 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3789 1063 1074 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3788 1339 1056 1063 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3787 1057 1058 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3786 1069 1059 1074 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3785 104 1059 1075 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3784 1074 1068 1062 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3783 1062 1075 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3782 1058 997 1061 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3781 1061 1081 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3780 1071 1057 1339 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3779 104 1057 1056 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3778 1339 1070 1060 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3777 1060 1056 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D3776 are shorted:
* D3776 104 104 D_lateral AREA=3.125E-016    $ (-592.5 608.499 -587.5 608.5)CMOSN3776 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3775 are shorted:
* D3775 88 88 D_lateral AREA=3.125E-016    $ (-603.5 533 -603.499 538)CMOSN3775 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3774 are shorted:
* D3774 88 88 D_lateral AREA=3.125E-016    $ (-654.5 622.499 -649.5 622.5)CMOSN3774 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3773 are shorted:
* D3773 88 88 D_lateral AREA=3.125E-016    $ (-608.5 622 -608.499 627)CMOSN3773 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3772 are shorted:
* D3772 88 88 D_lateral AREA=3.125E-016    $ (-648 578.499 -643 578.5)CMOSN3772 88 88 D_lateral AREA=3.125E-016    
M3771 88 1078 1072 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M3770 1073 1077 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3769 88 1081 1077 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3768 1068 1072 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3767 88 1072 1076 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3766 1076 1075 1074 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3765 88 997 1078 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3764 1070 1074 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3763 104 1078 1072 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M3762 1073 1077 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3761 1068 1072 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3760 104 1072 1069 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3758 1070 1074 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3757 104 1074 1071 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D3756 are shorted:
* D3756 88 88 D_lateral AREA=3.125E-016    $ (-780.5 578 -780.499 583)CMOSN3756 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3755 are shorted:
* D3755 104 104 D_lateral AREA=3.125E-016    $ (-723 608.499 -718 608.5)CMOSN3755 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3754 are shorted:
* D3754 88 88 D_lateral AREA=3.125E-016    $ (-780 622 -779.999 627)CMOSN3754 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3753 are shorted:
* D3753 104 104 D_lateral AREA=3.125E-016    $ (-716.5 564.499 -711.5 564.5)CMOSN3753 104 104 D_lateral AREA=3.125E-016    
M3752 1077 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3751 1078 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3750 88 1093 1084 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3749 1356 1345 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3748 88 1112 1345 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3746 1082 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3745 1077 1081 1082 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3744 1080 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3743 1080 997 1078 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3742 104 1093 1084 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3741 1345 1112 1079 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
* Pins of element D3739 are shorted:
* D3739 88 88 D_lateral AREA=3.125E-016    $ (-887.5 622.499 -882.5 622.5)CMOSN3739 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3738 are shorted:
* D3738 88 88 D_lateral AREA=3.125E-016    $ (-873 578 -872.999 583)CMOSN3738 88 88 D_lateral AREA=3.125E-016    
M3737 88 1093 1094 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3736 1094 1083 1086 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3735 1083 1102 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3734 88 1102 1092 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3733 1086 1084 1092 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3732 1091 1356 1110 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M3731 88 1346 1091 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M3730 1346 1344 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3729 88 1086 1345 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3728 88 1086 1344 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3727 1344 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3726 1101 1087 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3725 88 997 1087 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3724 1087 1112 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3723 1085 1093 1086 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3722 1086 1083 1090 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3721 104 1102 1085 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3720 1083 1102 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3719 1090 1084 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3718 104 1086 1079 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3717 1344 1086 1089 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3716 1089 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3715 1101 1087 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3714 1087 997 1088 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3713 1088 1112 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D3712 are shorted:
* D3712 104 104 D_lateral AREA=3.125E-016    $ (-956 608.499 -951 608.5)CMOSN3712 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3711 are shorted:
* D3711 88 88 D_lateral AREA=3.125E-016    $ (-967 533 -966.999 538)CMOSN3711 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3710 are shorted:
* D3710 88 88 D_lateral AREA=3.125E-016    $ (-917.5 578 -917.499 583)CMOSN3710 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3709 are shorted:
* D3709 88 88 D_lateral AREA=3.125E-016    $ (-972 622 -971.999 627)CMOSN3709 88 88 D_lateral AREA=3.125E-016    
M3708 1148 1355 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3707 1110 1113 1355 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M3706 88 1102 1096 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3705 88 1102 1109 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3704 1109 1095 1103 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3703 1095 1111 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3702 88 1111 1108 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3701 1103 1096 1108 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3700 88 1101 1099 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3699 88 1101 1107 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3698 1107 1098 1363 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3697 1098 1103 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3696 1106 1103 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3695 1363 1099 1106 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3694 1097 1102 1103 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3693 104 1102 1096 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3692 1103 1095 1105 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3691 104 1111 1097 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3690 1095 1111 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3689 1105 1096 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3688 1100 1101 1363 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3687 104 1101 1099 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3686 1363 1098 1104 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3685 104 1103 1100 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3684 1098 1103 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3683 1104 1099 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D3682 are shorted:
* D3682 88 88 D_lateral AREA=3.125E-016    $ (-1018 622.499 -1013 622.5)CMOSN3682 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3681 are shorted:
* D3681 104 104 D_lateral AREA=3.125E-016    $ (-1086.5 608.499 -1081.5 608.5)CMOSN3681 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3680 are shorted:
* D3680 88 88 D_lateral AREA=3.125E-016    $ (-1011.5 578.499 -1006.5 578.5)CMOSN3680 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3679 are shorted:
* D3679 104 104 D_lateral AREA=3.125E-016    $ (-1080 564.499 -1075 564.5)CMOSN3679 104 104 D_lateral AREA=3.125E-016    
M3678 88 1115 1111 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M3677 1113 1114 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3676 88 1112 1114 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3675 1114 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3674 88 997 1115 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3673 1115 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3672 104 1115 1111 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M3671 1113 1114 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3670 1114 1112 1117 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3669 1117 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3668 1115 997 1116 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3667 1116 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D3666 are shorted:
* D3666 88 88 D_lateral AREA=3.125E-016    $ (-1144 578 -1143.999 583)CMOSN3666 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3665 are shorted:
* D3665 88 88 D_lateral AREA=3.125E-016    $ (-1143.5 622 -1143.499 627)CMOSN3665 88 88 D_lateral AREA=3.125E-016    
M3664 88 1093 1129 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3663 88 1093 1119 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3662 1119 1124 1128 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3661 1367 1364 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3660 88 1148 1364 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3659 1364 1128 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3658 1120 1093 1128 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3657 104 1093 1129 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3655 1364 1148 1118 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3654 1118 1128 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D3653 are shorted:
* D3653 88 88 D_lateral AREA=3.125E-016    $ (-1259 622.499 -1254 622.5)CMOSN3653 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3652 are shorted:
* D3652 88 88 D_lateral AREA=3.125E-016    $ (-1244.5 578 -1244.499 583)CMOSN3652 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3651 are shorted:
* D3651 88 88 D_lateral AREA=3.125E-016    $ (-1289 578 -1288.999 583)CMOSN3651 88 88 D_lateral AREA=3.125E-016    
M3650 1124 1146 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3649 88 1146 1130 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3648 1128 1129 1130 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3647 1126 1367 1127 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M3646 88 1369 1126 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M3645 1127 1136 1379 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M3644 1369 1368 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3643 88 1128 1368 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3642 1368 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3641 1140 1121 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3639 88 997 1121 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3638 1121 1148 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3637 1138 1140 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M3636 1125 1124 1128 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=1.84375p PS=4.375u    
M3635 1124 1146 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3634 104 1146 1120 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3633 1125 1129 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3632 1368 1128 1123 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3631 1123 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3630 1140 1121 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3629 104 1146 1132 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3628 1121 997 1122 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3627 1122 1148 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3626 104 1140 1138 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D3625 are shorted:
* D3625 104 104 D_lateral AREA=3.125E-016    $ (-1327.5 608.499 -1322.5 608.5)CMOSN3625 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3624 are shorted:
* D3624 88 88 D_lateral AREA=3.125E-016    $ (-1338.5 533 -1338.499 538)CMOSN3624 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3623 are shorted:
* D3623 88 88 D_lateral AREA=3.125E-016    $ (-1389.5 622.499 -1384.5 622.5)CMOSN3623 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3622 are shorted:
* D3622 88 88 D_lateral AREA=3.125E-016    $ (-1343.5 622 -1343.499 627)CMOSN3622 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3621 are shorted:
* D3621 88 88 D_lateral AREA=3.125E-016    $ (-1383 578.499 -1378 578.5)CMOSN3621 88 88 D_lateral AREA=3.125E-016    
M3620 88 1150 1147 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M3619 1187 1379 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3618 1136 1149 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3617 1132 1146 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M3616 88 1146 1145 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3615 1145 1131 1137 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3614 1131 1147 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3613 88 1147 1144 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3612 1137 1132 1144 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3611 88 1140 1143 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3610 1143 1134 1385 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3609 1134 1137 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3608 1142 1137 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3607 1385 1138 1142 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3606 104 1150 1147 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M3605 1136 1149 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3604 1133 1146 1137 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3603 1137 1131 1141 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3602 104 1147 1133 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3601 1131 1147 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3600 1141 1132 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3599 1135 1140 1385 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3598 1385 1134 1139 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3597 104 1137 1135 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3596 1134 1137 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3595 1139 1138 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D3594 are shorted:
* D3594 104 104 D_lateral AREA=3.125E-016    $ (-1458 608.499 -1453 608.5)CMOSN3594 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3593 are shorted:
* D3593 104 104 D_lateral AREA=3.125E-016    $ (-1451.5 564.499 -1446.5 564.5)CMOSN3593 104 104 D_lateral AREA=3.125E-016    
M3592 88 1148 1149 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3591 1149 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3590 88 997 1150 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3589 1150 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3588 1149 1148 1152 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3587 1152 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3586 1150 997 1151 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3585 1151 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D3584 are shorted:
* D3584 88 88 D_lateral AREA=3.125E-016    $ (-1515.5 578 -1515.499 583)CMOSN3584 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3583 are shorted:
* D3583 88 88 D_lateral AREA=3.125E-016    $ (-1515 622 -1514.999 627)CMOSN3583 88 88 D_lateral AREA=3.125E-016    
M3582 88 1093 1154 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3581 88 1093 1161 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3580 1161 1153 1156 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3579 1153 1165 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3578 88 1165 1160 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3577 1156 1154 1160 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3576 1396 1390 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3575 1395 1391 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3574 88 1187 1391 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3573 1391 1156 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3572 88 1156 1390 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3571 1390 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3570 1155 1093 1156 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3569 104 1093 1154 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3568 1156 1153 1159 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3567 104 1165 1155 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3566 1153 1165 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3565 1159 1154 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3564 1391 1187 1158 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3563 1158 1156 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3562 1390 1156 1157 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3561 1157 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D3560 are shorted:
* D3560 88 88 D_lateral AREA=3.125E-016    $ (-1627 622.499 -1622 622.5)CMOSN3560 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3558 are shorted:
* D3558 88 88 D_lateral AREA=3.125E-016    $ (-1612.5 578 -1612.499 583)CMOSN3558 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3557 are shorted:
* D3557 88 88 D_lateral AREA=3.125E-016    $ (-1657 578 -1656.999 583)CMOSN3557 88 88 D_lateral AREA=3.125E-016    
M3556 1218 1402 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3555 1171 1395 1172 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M3554 88 1396 1171 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M3553 1172 1178 1402 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M3552 1163 1164 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3551 88 1165 1181 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3550 88 1165 1170 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3549 1170 1173 1180 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3548 88 997 1164 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3547 1164 1187 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3546 88 1163 1162 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3545 88 1163 1169 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3544 1169 1175 1408 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3542 1408 1162 1168 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3541 1163 1164 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3540 1174 1165 1180 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3539 104 1165 1181 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3538 1180 1173 1179 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3537 1164 997 1167 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3536 1167 1187 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3535 1176 1163 1408 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3534 104 1163 1162 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3533 1408 1175 1166 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3532 1166 1162 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D3531 are shorted:
* D3531 104 104 D_lateral AREA=3.125E-016    $ (-1695.5 608.499 -1690.5 608.5)CMOSN3531 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3530 are shorted:
* D3530 88 88 D_lateral AREA=3.125E-016    $ (-1706.5 533 -1706.499 538)CMOSN3530 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3529 are shorted:
* D3529 88 88 D_lateral AREA=3.125E-016    $ (-1757.5 622.499 -1752.5 622.5)CMOSN3529 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3528 are shorted:
* D3528 88 88 D_lateral AREA=3.125E-016    $ (-1711.5 622 -1711.499 627)CMOSN3528 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3527 are shorted:
* D3527 88 88 D_lateral AREA=3.125E-016    $ (-1751 578.499 -1746 578.5)CMOSN3527 88 88 D_lateral AREA=3.125E-016    
M3526 88 1184 1177 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M3525 1178 1183 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3523 1173 1177 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3522 88 1177 1182 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3521 1180 1181 1182 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3519 1175 1180 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3518 88 1180 1168 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3517 104 1184 1177 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M3516 1178 1183 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3515 1173 1177 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3514 104 1177 1174 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3513 1179 1181 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3512 1175 1180 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3511 104 1180 1176 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D3510 are shorted:
* D3510 88 88 D_lateral AREA=3.125E-016    $ (-1883.5 578 -1883.499 583)CMOSN3510 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3509 are shorted:
* D3509 104 104 D_lateral AREA=3.125E-016    $ (-1826 608.499 -1821 608.5)CMOSN3509 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3508 are shorted:
* D3508 88 88 D_lateral AREA=3.125E-016    $ (-1883 622 -1882.999 627)CMOSN3508 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3507 are shorted:
* D3507 104 104 D_lateral AREA=3.125E-016    $ (-1819.5 564.499 -1814.5 564.5)CMOSN3507 104 104 D_lateral AREA=3.125E-016    
M3506 1422 1195 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3505 88 1218 1195 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3504 1183 1187 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3503 1183 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3502 1184 997 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3501 1184 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3499 1195 1218 1193 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3498 1183 1187 1186 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3497 1186 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3496 1184 997 1185 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3495 1185 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D3494 are shorted:
* D3494 88 88 D_lateral AREA=3.125E-016    $ (-1991 622.499 -1986 622.5)CMOSN3494 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3493 are shorted:
* D3493 88 88 D_lateral AREA=3.125E-016    $ (-1976.5 578 -1976.499 583)CMOSN3493 88 88 D_lateral AREA=3.125E-016    
M3492 88 1093 1189 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3491 88 1093 1198 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3490 1198 1188 1191 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3489 1188 1206 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3488 88 1206 1197 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3487 1191 1189 1197 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3485 88 1414 1196 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M3484 1414 1413 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3483 1195 1191 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3482 88 1191 1413 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3481 1413 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3480 1205 1213 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3479 88 997 1213 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3478 1190 1093 1191 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3477 1189 1093 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3476 1191 1188 1194 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3475 104 1206 1190 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3474 1188 1206 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3473 1194 1189 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3472 1193 1191 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3471 1413 1191 1192 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3470 1192 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3469 1205 1213 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3468 1213 997 1209 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
* Pins of element D3467 are shorted:
* D3467 104 104 D_lateral AREA=3.125E-016    $ (-2059.5 608.499 -2054.5 608.5)CMOSN3467 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3466 are shorted:
* D3466 88 88 D_lateral AREA=3.125E-016    $ (-2070.5 533 -2070.499 538)CMOSN3466 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3465 are shorted:
* D3465 88 88 D_lateral AREA=3.125E-016    $ (-2021 578 -2020.999 583)CMOSN3465 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3464 are shorted:
* D3464 88 88 D_lateral AREA=3.125E-016    $ (-2075.5 622 -2075.499 627)CMOSN3464 88 88 D_lateral AREA=3.125E-016    
M3463 1254 1421 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3462 1216 1422 1196 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.125p PS=3.75u    
M3461 1216 1219 1421 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M3460 88 1206 1200 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3459 88 1206 1215 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3458 1215 1199 1207 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3457 1199 1217 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3456 88 1217 1214 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3455 1207 1200 1214 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3454 1213 1218 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3453 88 1205 1203 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3452 88 1205 1212 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3451 1212 1202 1431 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3450 1202 1207 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3449 1211 1207 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3448 1431 1203 1211 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3447 1201 1206 1207 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3446 104 1206 1200 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3445 1207 1199 1210 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3444 104 1217 1201 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3443 1199 1217 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3442 1210 1200 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3441 1209 1218 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3440 1204 1205 1431 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3439 104 1205 1203 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3438 1431 1202 1208 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3437 104 1207 1204 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3436 1202 1207 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3435 1208 1203 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D3434 are shorted:
* D3434 88 88 D_lateral AREA=3.125E-016    $ (-2121.5 622.499 -2116.5 622.5)CMOSN3434 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3433 are shorted:
* D3433 104 104 D_lateral AREA=3.125E-016    $ (-2190 608.499 -2185 608.5)CMOSN3433 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3432 are shorted:
* D3432 88 88 D_lateral AREA=3.125E-016    $ (-2115 578.499 -2110 578.5)CMOSN3432 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3431 are shorted:
* D3431 104 104 D_lateral AREA=3.125E-016    $ (-2183.5 564.499 -2178.5 564.5)CMOSN3431 104 104 D_lateral AREA=3.125E-016    
M3430 88 1221 1217 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M3429 1219 1220 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3428 88 1218 1220 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3427 1220 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3426 88 997 1221 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3425 1221 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3424 104 1221 1217 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M3423 1219 1220 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3422 1220 1218 1223 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3421 1223 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3420 1221 997 1222 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3419 1222 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D3418 are shorted:
* D3418 88 88 D_lateral AREA=3.125E-016    $ (-2247.5 578 -2247.499 583)CMOSN3418 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3417 are shorted:
* D3417 88 88 D_lateral AREA=3.125E-016    $ (-2247 622 -2246.999 627)CMOSN3417 88 88 D_lateral AREA=3.125E-016    
M3416 88 1093 1235 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3415 88 1093 1225 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3414 1225 1230 1234 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3413 1435 1432 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3412 88 1254 1432 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3411 1432 1234 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3410 1226 1093 1234 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3409 104 1093 1235 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3408 1432 1254 1224 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3407 1224 1234 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D3406 are shorted:
* D3406 88 88 D_lateral AREA=3.125E-016    $ (-2361.5 622.499 -2356.5 622.5)CMOSN3406 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3405 are shorted:
* D3405 88 88 D_lateral AREA=3.125E-016    $ (-2347 578 -2346.999 583)CMOSN3405 88 88 D_lateral AREA=3.125E-016    
M3404 1230 1241 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3403 88 1241 1236 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3402 1234 1235 1236 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3401 1232 1435 1233 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M3400 88 1437 1232 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M3399 1233 1244 1447 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M3398 1437 1436 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3397 88 1234 1436 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3396 1436 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3395 1247 1227 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3394 88 997 1227 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3393 1227 1254 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3392 1237 1247 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M3391 1234 1230 1231 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3390 104 1241 1226 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3389 1230 1241 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3388 1231 1235 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3387 1436 1234 1229 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3386 1229 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3385 1247 1227 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3383 1227 997 1228 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3382 1228 1254 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3381 104 1247 1237 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D3380 are shorted:
* D3380 104 104 D_lateral AREA=3.125E-016    $ (-2430 608.499 -2425 608.5)CMOSN3380 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3379 are shorted:
* D3379 88 88 D_lateral AREA=3.125E-016    $ (-2441 533 -2440.999 538)CMOSN3379 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3378 are shorted:
* D3378 88 88 D_lateral AREA=3.125E-016    $ (-2391.5 578 -2391.499 583)CMOSN3378 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3376 are shorted:
* D3376 88 88 D_lateral AREA=3.125E-016    $ (-2446 622 -2445.999 627)CMOSN3376 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3375 are shorted:
* D3375 88 88 D_lateral AREA=3.125E-016    $ (-2485.5 578.499 -2480.5 578.5)CMOSN3375 88 88 D_lateral AREA=3.125E-016    
M3374 88 1256 1253 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M3373 1475 1447 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3372 1244 1255 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M3371 88 1241 1239 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3370 88 1241 1252 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3369 1252 1238 1245 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3368 1238 1253 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3367 88 1253 1251 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3366 1245 1239 1251 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3365 88 1247 1250 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3364 1250 1242 1452 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3363 1242 1245 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3362 1249 1245 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3361 1452 1237 1249 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3360 104 1256 1253 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M3359 1244 1255 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3358 1240 1241 1245 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3357 1239 1241 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3356 1245 1238 1248 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3355 104 1253 1240 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3354 1238 1253 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3353 1248 1239 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3352 1243 1247 1452 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3351 1452 1242 1246 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3350 104 1245 1243 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3349 1242 1245 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3348 1246 1237 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D3347 are shorted:
* D3347 88 88 D_lateral AREA=3.125E-016    $ (-2492 622.499 -2487 622.5)CMOSN3347 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3346 are shorted:
* D3346 104 104 D_lateral AREA=3.125E-016    $ (-2560.5 608.499 -2555.5 608.5)CMOSN3346 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3345 are shorted:
* D3345 104 104 D_lateral AREA=3.125E-016    $ (-2554 564.499 -2549 564.5)CMOSN3345 104 104 D_lateral AREA=3.125E-016    
M3344 88 1254 1255 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3343 1255 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3342 88 997 1256 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3341 1256 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3340 1255 1254 1258 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3339 1258 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3338 1256 997 1257 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3337 1257 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D3336 are shorted:
* D3336 88 88 D_lateral AREA=3.125E-016    $ (-2618 578 -2617.999 583)CMOSN3336 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3335 are shorted:
* D3335 88 88 D_lateral AREA=3.125E-016    $ (-2617.5 622 -2617.499 627)CMOSN3335 88 88 D_lateral AREA=3.125E-016    
M3334 88 1093 1468 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3333 88 1093 1264 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3332 1093 1259 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M3331 997 1260 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M3330 1093 1259 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3329 997 1260 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D3328 are shorted:
* D3328 88 88 D_lateral AREA=3.125E-016    $ (-2870.5 531.999 -2865.5 532)CMOSN3328 88 88 D_lateral AREA=3.125E-016    
M3327 1470 1469 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3326 1265 1469 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3325 1264 1470 1481 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3324 1481 1468 1265 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3323 1469 1476 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M3322 88 976 1259 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3321 1259 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3320 1263 491 88 88 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M3319 1260 1261 1263 88 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M3318 1261 1271 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M3317 88 1269 1271 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3316 994 1266 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M3315 1259 976 1262 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3314 1262 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3313 1260 491 104 104 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M3312 104 1261 1260 104 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M3311 1261 1271 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3309 994 1266 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D3308 are shorted:
* D3308 88 88 D_lateral AREA=3.125E-016    $ (-2893.5 576.5 -2893.499 581.5)CMOSN3308 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3307 are shorted:
* D3307 88 88 D_lateral AREA=3.125E-016    $ (-2977.5 576.5 -2977.499 581.5)CMOSN3307 88 88 D_lateral AREA=3.125E-016    
M3306 88 1475 1476 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3305 1476 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3304 1271 1267 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3303 1267 491 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M3302 88 1269 1266 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3301 1266 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3300 1270 1267 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3299 1270 1269 1271 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3298 1267 491 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3297 1266 1269 1268 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3296 1268 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D3295 are shorted:
* D3295 88 88 D_lateral AREA=3.125E-016    $ (-2998.5 531.5 -2998.499 536.5)CMOSN3295 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3294 are shorted:
* D3294 88 88 D_lateral AREA=3.125E-016    $ (-3006.5 622 -3006.499 627)CMOSN3294 88 88 D_lateral AREA=3.125E-016    
M3292 88 1349 1273 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3291 88 1349 1280 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3290 1280 1272 1489 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3289 1272 1284 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3288 1279 1284 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3287 1489 1273 1279 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3286 88 1287 1498 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3285 1274 1349 1489 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3284 104 1349 1273 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3283 1489 1272 1278 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3282 104 1284 1274 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3281 1272 1284 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3280 1278 1273 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3279 104 1277 1285 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M3278 1277 1275 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3277 104 1276 1286 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D3276 are shorted:
* D3276 88 88 D_lateral AREA=3.125E-016    $ (203.5 459.999 208.5 460)CMOSN3276 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3275 are shorted:
* D3275 104 104 D_lateral AREA=3.125E-016    $ (135 445.999 140 446)CMOSN3275 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3274 are shorted:
* D3274 88 88 D_lateral AREA=3.125E-016    $ (119 459.5 119.001 464.5)CMOSN3274 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3273 are shorted:
* D3273 104 104 D_lateral AREA=3.125E-016    $ (125.999 516 126 521)CMOSN3273 104 104 D_lateral AREA=3.125E-016    
M3272 88 1284 1282 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3271 88 1284 1291 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3270 1291 1281 1499 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3269 1281 1292 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3268 1290 1292 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3267 1499 1282 1290 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3266 1498 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3265 1283 1284 1499 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3264 104 1284 1282 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3263 1499 1281 1289 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3262 104 1292 1283 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3261 1281 1292 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3260 1289 1282 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3259 1288 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3258 1498 1287 1288 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3257 1042 1285 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3256 1285 1286 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M3255 104 1007 1285 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
* Pins of element D3254 are shorted:
* D3254 88 88 D_lateral AREA=3.125E-016    $ (73 459.999 78 460)CMOSN3254 88 88 D_lateral AREA=3.125E-016    
M3252 88 1293 1292 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M3251 88 1287 1293 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3250 1293 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3249 104 1293 1292 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M3248 1293 1287 1294 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3247 1294 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D3246 are shorted:
* D3246 104 104 D_lateral AREA=3.125E-016    $ (4.5 445.999 9.5 446)CMOSN3246 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3245 are shorted:
* D3245 88 88 D_lateral AREA=3.125E-016    $ (-52.5 459.5 -52.499 464.5)CMOSN3245 88 88 D_lateral AREA=3.125E-016    
M3244 88 1349 1306 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3243 88 1349 1297 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3242 1297 1303 1305 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3241 1298 1349 1305 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3240 104 1349 1306 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3238 1299 1296 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D3237 are shorted:
* D3237 88 88 D_lateral AREA=3.125E-016    $ (-160 459.999 -155 460)CMOSN3237 88 88 D_lateral AREA=3.125E-016    
M3236 1303 1295 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3235 1307 1295 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3234 1305 1306 1307 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3233 88 1287 1513 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3232 1513 1528 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3231 1304 1303 1305 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=1.84375p PS=4.375u    
M3230 1303 1295 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3229 104 1295 1298 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3228 1304 1306 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3227 104 1295 1309 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3226 1513 1287 1302 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3225 1302 1528 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3224 1311 1299 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M3223 104 1031 1311 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M3222 104 1301 1311 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M3221 1301 1300 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D3220 are shorted:
* D3220 104 104 D_lateral AREA=3.125E-016    $ (-228.5 445.999 -223.5 446)CMOSN3220 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3219 are shorted:
* D3219 88 88 D_lateral AREA=3.125E-016    $ (-290.5 459.999 -285.5 460)CMOSN3219 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3218 are shorted:
* D3218 88 88 D_lateral AREA=3.125E-016    $ (-244.5 459.5 -244.499 464.5)CMOSN3218 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3217 are shorted:
* D3217 104 104 D_lateral AREA=3.125E-016    $ (-237.501 516 -237.5 521)CMOSN3217 104 104 D_lateral AREA=3.125E-016    
M3216 88 1315 1316 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M3215 88 1295 1309 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3214 88 1295 1314 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3213 1314 1308 1522 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3212 1308 1316 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3211 1313 1316 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3210 1522 1309 1313 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3209 104 1315 1316 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M3208 1310 1295 1522 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3207 1522 1308 1312 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3206 104 1316 1310 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3205 1308 1316 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3204 1312 1309 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3203 1081 1311 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D3202 are shorted:
* D3202 104 104 D_lateral AREA=3.125E-016    $ (-359 445.999 -354 446)CMOSN3202 104 104 D_lateral AREA=3.125E-016    
M3201 88 1287 1315 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3200 1315 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3199 1315 1287 1318 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3198 1318 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D3197 are shorted:
* D3197 88 88 D_lateral AREA=3.125E-016    $ (-416 459.5 -415.999 464.5)CMOSN3197 88 88 D_lateral AREA=3.125E-016    
M3196 88 1349 1320 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3195 88 1349 1326 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3194 1326 1319 1532 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3193 1319 1317 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3192 1325 1317 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3191 1532 1320 1325 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3190 1321 1349 1532 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3189 104 1349 1320 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3188 1532 1319 1324 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3187 104 1317 1321 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3186 1319 1317 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3185 1324 1320 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3184 1329 1322 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3183 1328 1323 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D3182 are shorted:
* D3182 88 88 D_lateral AREA=3.125E-016    $ (-524.5 459.999 -519.5 460)CMOSN3182 88 88 D_lateral AREA=3.125E-016    
M3180 88 1317 1336 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3179 88 1317 1332 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3178 1332 1333 1549 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3176 88 1287 1539 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3175 1539 1552 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3174 1334 1317 1549 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3173 104 1317 1336 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3172 1549 1333 1331 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3170 1539 1287 1330 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3169 1330 1552 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3168 1112 1327 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3167 1327 1328 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M3166 104 1073 1327 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M3165 104 1329 1327 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
* Pins of element D3164 are shorted:
* D3164 104 104 D_lateral AREA=3.125E-016    $ (-593 445.999 -588 446)CMOSN3164 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3163 are shorted:
* D3163 88 88 D_lateral AREA=3.125E-016    $ (-655 459.999 -650 460)CMOSN3163 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3162 are shorted:
* D3162 88 88 D_lateral AREA=3.125E-016    $ (-609 459.5 -608.999 464.5)CMOSN3162 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3161 are shorted:
* D3161 104 104 D_lateral AREA=3.125E-016    $ (-602.001 516 -602 521)CMOSN3161 104 104 D_lateral AREA=3.125E-016    
M3160 88 1338 1335 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M3159 1333 1335 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3158 1337 1335 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3157 1337 1336 1549 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3156 88 1287 1338 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3155 104 1338 1335 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M3154 1333 1335 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3153 104 1335 1334 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3152 104 1336 1331 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=187.5f PS=1.25u    
* Pins of element D3151 are shorted:
* D3151 104 104 D_lateral AREA=3.125E-016    $ (-723.5 445.999 -718.5 446)CMOSN3151 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3150 are shorted:
* D3150 88 88 D_lateral AREA=3.125E-016    $ (-780.5 459.5 -780.499 464.5)CMOSN3150 88 88 D_lateral AREA=3.125E-016    
M3149 1338 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3148 1342 1349 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M3147 1340 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3146 1338 1287 1340 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3145 104 1349 1342 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3144 1356 1345 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D3143 are shorted:
* D3143 88 88 D_lateral AREA=3.125E-016    $ (-888 459.999 -883 460)CMOSN3143 88 88 D_lateral AREA=3.125E-016    
M3142 88 1349 1351 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3141 1351 1341 1557 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3140 1341 1339 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3139 1350 1339 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3138 1557 1342 1350 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3137 88 1287 1558 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3135 1343 1349 1557 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3134 1557 1341 1348 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3133 104 1339 1343 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3132 1341 1339 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3131 1348 1342 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3130 1558 1287 1347 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3127 104 1346 1355 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M3126 1346 1344 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D3125 are shorted:
* D3125 104 104 D_lateral AREA=3.125E-016    $ (-956.5 445.999 -951.5 446)CMOSN3125 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3124 are shorted:
* D3124 88 88 D_lateral AREA=3.125E-016    $ (-972.5 459.5 -972.499 464.5)CMOSN3124 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3123 are shorted:
* D3123 104 104 D_lateral AREA=3.125E-016    $ (-965.501 516 -965.5 521)CMOSN3123 104 104 D_lateral AREA=3.125E-016    
M3122 88 1339 1353 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3121 88 1339 1359 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3120 1359 1352 1566 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3119 1352 1361 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3118 1358 1361 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3117 1566 1353 1358 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3116 88 1574 1558 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3115 1354 1339 1566 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3114 104 1339 1353 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3113 1566 1352 1357 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3112 104 1361 1354 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3111 1352 1361 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3110 1357 1353 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3109 104 1574 1347 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3108 1148 1355 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3107 104 1113 1355 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M3106 104 1356 1355 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=1.15625p PS=3.5u    
* Pins of element D3105 are shorted:
* D3105 88 88 D_lateral AREA=3.125E-016    $ (-1018.5 459.999 -1013.5 460)CMOSN3105 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3104 are shorted:
* D3104 104 104 D_lateral AREA=3.125E-016    $ (-1087 445.999 -1082 446)CMOSN3104 104 104 D_lateral AREA=3.125E-016    
M3103 88 1360 1361 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M3102 88 1287 1360 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3101 1360 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3100 104 1360 1361 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M3099 1360 1287 1362 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3098 1362 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D3097 are shorted:
* D3097 88 88 D_lateral AREA=3.125E-016    $ (-1144 459.5 -1143.999 464.5)CMOSN3097 88 88 D_lateral AREA=3.125E-016    
M3096 88 1349 1374 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3095 88 1349 1365 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3094 1365 1371 1373 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3093 1366 1349 1373 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3092 104 1349 1374 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3090 1367 1364 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D3089 are shorted:
* D3089 88 88 D_lateral AREA=3.125E-016    $ (-1259.5 459.999 -1254.5 460)CMOSN3089 88 88 D_lateral AREA=3.125E-016    
M3088 1371 1363 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3087 1375 1363 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3086 1373 1374 1375 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3084 88 1287 1581 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3083 1581 1596 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3082 1372 1371 1373 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=1.84375p PS=4.375u    
M3081 1371 1363 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3080 104 1363 1366 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3079 1372 1374 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3078 104 1363 1377 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3077 1581 1287 1370 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3076 1370 1596 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3075 1379 1367 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M3074 104 1136 1379 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M3073 104 1369 1379 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M3072 1369 1368 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D3071 are shorted:
* D3071 104 104 D_lateral AREA=3.125E-016    $ (-1328 445.999 -1323 446)CMOSN3071 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3070 are shorted:
* D3070 88 88 D_lateral AREA=3.125E-016    $ (-1390 459.999 -1385 460)CMOSN3070 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3069 are shorted:
* D3069 88 88 D_lateral AREA=3.125E-016    $ (-1344 459.5 -1343.999 464.5)CMOSN3069 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3068 are shorted:
* D3068 104 104 D_lateral AREA=3.125E-016    $ (-1337.001 516 -1337 521)CMOSN3068 104 104 D_lateral AREA=3.125E-016    
M3067 88 1383 1384 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M3066 1377 1363 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M3065 88 1363 1382 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3064 1382 1376 1590 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3063 1376 1384 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3062 1381 1384 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3061 1590 1377 1381 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3060 104 1383 1384 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M3059 1378 1363 1590 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3058 1590 1376 1380 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3057 104 1384 1378 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3056 1376 1384 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3055 1380 1377 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3054 1187 1379 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D3053 are shorted:
* D3053 104 104 D_lateral AREA=3.125E-016    $ (-1458.5 445.999 -1453.5 446)CMOSN3053 104 104 D_lateral AREA=3.125E-016    
M3052 88 1287 1383 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3051 1383 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3050 1383 1287 1386 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3049 1386 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D3048 are shorted:
* D3048 88 88 D_lateral AREA=3.125E-016    $ (-1515.5 459.5 -1515.499 464.5)CMOSN3048 88 88 D_lateral AREA=3.125E-016    
M3047 88 1349 1388 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3046 88 1349 1394 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3045 1394 1387 1600 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3044 1387 1385 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3043 1393 1385 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3042 1600 1388 1393 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3041 1389 1349 1600 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3040 104 1349 1388 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3039 1600 1387 1392 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3038 104 1385 1389 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3037 1387 1385 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3036 1392 1388 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M3035 1396 1390 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3034 1395 1391 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D3033 are shorted:
* D3033 88 88 D_lateral AREA=3.125E-016    $ (-1627.5 459.999 -1622.5 460)CMOSN3033 88 88 D_lateral AREA=3.125E-016    
M3031 88 1385 1405 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M3030 88 1385 1398 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M3029 1398 1399 1404 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M3028 88 1287 1607 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3027 1607 1619 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3026 1400 1385 1404 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M3025 104 1385 1405 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3024 1404 1399 1403 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M3023 1607 1287 1397 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3022 1397 1619 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3021 1218 1402 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M3020 1402 1395 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M3019 104 1178 1402 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M3018 104 1396 1402 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
* Pins of element D3017 are shorted:
* D3017 104 104 D_lateral AREA=3.125E-016    $ (-1696 445.999 -1691 446)CMOSN3017 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3016 are shorted:
* D3016 88 88 D_lateral AREA=3.125E-016    $ (-1758 459.999 -1753 460)CMOSN3016 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3015 are shorted:
* D3015 88 88 D_lateral AREA=3.125E-016    $ (-1712 459.5 -1711.999 464.5)CMOSN3015 88 88 D_lateral AREA=3.125E-016    
* Pins of element D3014 are shorted:
* D3014 104 104 D_lateral AREA=3.125E-016    $ (-1705.001 516 -1705 521)CMOSN3014 104 104 D_lateral AREA=3.125E-016    
M3013 88 1407 1401 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M3012 1399 1401 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3011 1406 1401 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3010 1404 1405 1406 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M3008 104 1407 1401 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M3007 1399 1401 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M3006 104 1401 1400 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3005 1403 1405 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D3004 are shorted:
* D3004 104 104 D_lateral AREA=3.125E-016    $ (-1826.5 445.999 -1821.5 446)CMOSN3004 104 104 D_lateral AREA=3.125E-016    
* Pins of element D3003 are shorted:
* D3003 88 88 D_lateral AREA=3.125E-016    $ (-1883.5 459.5 -1883.499 464.5)CMOSN3003 88 88 D_lateral AREA=3.125E-016    
M3002 1407 1287 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3001 1407 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2999 1407 1287 1409 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2998 1409 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2997 1422 1195 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2995 88 1349 1411 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2994 88 1349 1417 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2993 1417 1410 1622 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2992 1410 1408 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2991 1416 1408 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2990 1622 1411 1416 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2989 88 1287 1425 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2988 1412 1349 1622 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2987 1411 1349 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2986 1622 1410 1415 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2985 104 1408 1412 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2984 1410 1408 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2983 1415 1411 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M2982 1425 1287 1423 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2980 104 1414 1421 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M2979 1414 1413 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D2978 are shorted:
* D2978 88 88 D_lateral AREA=3.125E-016    $ (-1991.5 459.999 -1986.5 460)CMOSN2978 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2977 are shorted:
* D2977 104 104 D_lateral AREA=3.125E-016    $ (-2060 445.999 -2055 446)CMOSN2977 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2976 are shorted:
* D2976 88 88 D_lateral AREA=3.125E-016    $ (-2076 459.5 -2075.999 464.5)CMOSN2976 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2975 are shorted:
* D2975 104 104 D_lateral AREA=3.125E-016    $ (-2069.001 516 -2069 521)CMOSN2975 104 104 D_lateral AREA=3.125E-016    
M2974 88 1408 1419 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2973 88 1408 1427 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2972 1427 1418 1632 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2971 1418 1429 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2970 1426 1429 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2969 1632 1419 1426 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2968 1425 1640 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2967 1420 1408 1632 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2966 104 1408 1419 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2965 1632 1418 1424 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2964 104 1429 1420 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2963 1418 1429 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2962 1424 1419 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M2961 1423 1640 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2960 1254 1421 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2959 104 1422 1421 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=1.15625p PS=3.5u    
M2958 104 1219 1421 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
* Pins of element D2957 are shorted:
* D2957 88 88 D_lateral AREA=3.125E-016    $ (-2122 459.999 -2117 460)CMOSN2957 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2956 are shorted:
* D2956 104 104 D_lateral AREA=3.125E-016    $ (-2190.5 445.999 -2185.5 446)CMOSN2956 104 104 D_lateral AREA=3.125E-016    
M2955 88 1428 1429 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2954 88 1287 1428 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2953 1428 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2952 104 1428 1429 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2951 1428 1287 1430 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2950 1430 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2949 are shorted:
* D2949 88 88 D_lateral AREA=3.125E-016    $ (-2247.5 459.5 -2247.499 464.5)CMOSN2949 88 88 D_lateral AREA=3.125E-016    
M2948 88 1349 1442 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2947 88 1349 1433 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2946 1433 1439 1441 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2945 1434 1349 1441 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2944 104 1349 1442 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2943 1435 1432 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D2942 are shorted:
* D2942 88 88 D_lateral AREA=3.125E-016    $ (-2362 459.999 -2357 460)CMOSN2942 88 88 D_lateral AREA=3.125E-016    
M2941 1439 1431 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2940 1443 1431 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2939 1441 1442 1443 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2938 88 1287 1647 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2937 1647 1662 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2936 1441 1439 1440 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2935 104 1431 1434 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2934 1439 1431 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2933 1440 1442 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M2931 1647 1287 1438 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2930 1438 1662 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2929 1447 1435 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M2928 104 1244 1447 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M2927 104 1437 1447 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M2926 1437 1436 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D2925 are shorted:
* D2925 104 104 D_lateral AREA=3.125E-016    $ (-2430.5 445.999 -2425.5 446)CMOSN2925 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2923 are shorted:
* D2923 88 88 D_lateral AREA=3.125E-016    $ (-2446.5 459.5 -2446.499 464.5)CMOSN2923 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2922 are shorted:
* D2922 104 104 D_lateral AREA=3.125E-016    $ (-2439.501 516 -2439.5 521)CMOSN2922 104 104 D_lateral AREA=3.125E-016    
M2920 88 1431 1445 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2919 88 1431 1450 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2918 1450 1444 1656 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2917 1444 1451 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2916 1449 1451 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2915 1656 1445 1449 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2913 1446 1431 1656 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2912 1445 1431 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2911 1656 1444 1448 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2910 104 1451 1446 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2909 1444 1451 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2908 1448 1445 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M2907 1475 1447 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D2906 are shorted:
* D2906 88 88 D_lateral AREA=3.125E-016    $ (-2492.5 459.999 -2487.5 460)CMOSN2906 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2905 are shorted:
* D2905 104 104 D_lateral AREA=3.125E-016    $ (-2561 445.999 -2556 446)CMOSN2905 104 104 D_lateral AREA=3.125E-016    
M2904 1451 1454 88 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2903 88 1287 1454 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2902 1454 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2901 1451 1454 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.90625p PS=5.75u    
M2900 1454 1287 1453 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2899 1453 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2898 are shorted:
* D2898 88 88 D_lateral AREA=3.125E-016    $ (-2618 459.5 -2617.999 464.5)CMOSN2898 88 88 D_lateral AREA=3.125E-016    
M2897 88 1349 1456 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2896 88 1349 1460 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2895 1460 1455 1666 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2894 1455 1452 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2893 1459 1452 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2892 1666 1456 1459 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2891 1457 1349 1666 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2890 104 1349 1456 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2889 1666 1455 1458 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2888 104 1452 1457 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2886 1458 1456 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D2885 are shorted:
* D2885 88 88 D_lateral AREA=3.125E-016    $ (-2729 459.999 -2724 460)CMOSN2885 88 88 D_lateral AREA=3.125E-016    
M2884 88 1452 1473 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2883 88 1452 1462 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2882 1462 1466 1472 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2881 88 1287 1673 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2880 1673 1683 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2879 1463 1093 1481 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2878 104 1093 1468 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2877 104 1452 1455 104 CMOSN L=500n W=750n AD=2.21875p PD=6.25u AS=1.75p PS=5.5u    
M2876 1464 1452 1472 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2875 104 1452 1473 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2873 1673 1287 1461 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2872 1461 1683 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2871 are shorted:
* D2871 104 104 D_lateral AREA=3.125E-016    $ (-2797.5 445.999 -2792.5 446)CMOSN2871 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2870 are shorted:
* D2870 88 88 D_lateral AREA=3.125E-016    $ (-2859.5 459.999 -2854.5 460)CMOSN2870 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2869 are shorted:
* D2869 88 88 D_lateral AREA=3.125E-016    $ (-2813.5 459.5 -2813.499 464.5)CMOSN2869 88 88 D_lateral AREA=3.125E-016    
M2868 88 1477 1465 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2867 1466 1465 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2866 1474 1465 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2865 1472 1473 1474 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2863 1481 1470 1471 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2862 104 1469 1463 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2861 1470 1469 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2860 1471 1468 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M2859 1469 1476 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2858 104 1477 1465 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2857 1467 1466 1472 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=1.84375p PS=4.375u    
M2856 1466 1465 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2855 104 1465 1464 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2854 1467 1473 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D2853 are shorted:
* D2853 104 104 D_lateral AREA=3.125E-016    $ (-2939 517.999 -2934 518)CMOSN2853 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2852 are shorted:
* D2852 104 104 D_lateral AREA=3.125E-016    $ (-2928 445.999 -2923 446)CMOSN2852 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2851 are shorted:
* D2851 88 88 D_lateral AREA=3.125E-016    $ (-2985 459.5 -2984.999 464.5)CMOSN2851 88 88 D_lateral AREA=3.125E-016    
M2850 1477 1287 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2849 1477 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2848 1476 1475 1479 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2847 1479 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2846 1477 1287 1478 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2845 1478 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2844 1287 1480 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M2843 1287 1480 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2842 1482 491 88 88 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M2841 1480 1698 1482 88 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M2840 1284 1483 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M2839 88 1484 1483 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2838 1480 491 104 104 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M2837 104 1698 1480 104 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M2836 1284 1483 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D2835 are shorted:
* D2835 88 88 D_lateral AREA=3.125E-016    $ (-3381 459.5 -3380.999 464.5)CMOSN2835 88 88 D_lateral AREA=3.125E-016    
M2834 1483 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2833 1485 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2832 1483 1484 1485 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2830 88 104 1488 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
* Pins of element D2828 are shorted:
* D2828 88 88 D_lateral AREA=3.125E-016    $ (218 415.5 218.001 420.5)CMOSN2828 88 88 D_lateral AREA=3.125E-016    
M2827 88 1486 1503 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M2826 1486 1487 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2825 88 1488 1497 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2824 1488 1489 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2823 88 1489 1487 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2822 1487 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2821 1495 1498 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2820 104 1486 1496 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M2819 1486 1487 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2818 104 1488 1497 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2817 1488 104 1491 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2816 1491 1489 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2815 1487 1489 1490 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2814 1490 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2813 1495 1498 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D2812 are shorted:
* D2812 88 88 D_lateral AREA=3.125E-016    $ (124 370.5 124.001 375.5)CMOSN2812 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2811 are shorted:
* D2811 104 104 D_lateral AREA=3.125E-016    $ (125.499 353.5 125.5 358.5)CMOSN2811 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2810 are shorted:
* D2810 88 88 D_lateral AREA=3.125E-016    $ (173.5 415.5 173.501 420.5)CMOSN2810 88 88 D_lateral AREA=3.125E-016    
M2809 1528 1496 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2808 1503 1497 1504 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M2807 1504 1505 1496 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M2806 88 1495 1493 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2805 88 1495 1502 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2804 1502 1492 1747 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2803 1492 1499 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2802 1501 1499 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2801 1747 1493 1501 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2800 1528 1496 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2799 1496 1497 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M2798 104 1505 1496 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M2797 1494 1495 1747 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2796 104 1495 1493 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2795 1747 1492 1500 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2794 104 1499 1494 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2793 1492 1499 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2792 1500 1493 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D2791 are shorted:
* D2791 88 88 D_lateral AREA=3.125E-016    $ (79.5 415.999 84.5 416)CMOSN2791 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2790 are shorted:
* D2790 104 104 D_lateral AREA=3.125E-016    $ (11 401.999 16 402)CMOSN2790 104 104 D_lateral AREA=3.125E-016    
M2789 1505 1506 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2788 88 104 1506 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2787 1506 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2786 1505 1506 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2785 1506 104 1507 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2784 1507 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2783 are shorted:
* D2783 88 88 D_lateral AREA=3.125E-016    $ (-53 415.5 -52.999 420.5)CMOSN2783 88 88 D_lateral AREA=3.125E-016    
M2782 1510 1508 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2781 88 1528 1508 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2780 1508 1305 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2779 1510 1508 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2778 1508 1528 1509 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2777 1509 1305 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2776 are shorted:
* D2776 88 88 D_lateral AREA=3.125E-016    $ (-145.5 415.5 -145.499 420.5)CMOSN2776 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2775 are shorted:
* D2775 88 88 D_lateral AREA=3.125E-016    $ (-190 415.5 -189.999 420.5)CMOSN2775 88 88 D_lateral AREA=3.125E-016    
M2774 1515 1510 1516 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M2773 88 1511 1515 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M2772 1516 1520 1521 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M2771 1511 1512 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2770 88 1305 1512 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2769 1512 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2768 1524 1513 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2767 1518 1524 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M2766 1521 1510 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M2765 104 1511 1521 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M2764 104 1520 1521 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M2763 1511 1512 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2762 1512 1305 1514 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2761 1514 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2760 1524 1513 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2759 104 1524 1518 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D2758 are shorted:
* D2758 104 104 D_lateral AREA=3.125E-016    $ (-238.001 353.5 -238 358.5)CMOSN2758 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2757 are shorted:
* D2757 88 88 D_lateral AREA=3.125E-016    $ (-239.5 370.5 -239.499 375.5)CMOSN2757 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2756 are shorted:
* D2756 88 88 D_lateral AREA=3.125E-016    $ (-284 415.999 -279 416)CMOSN2756 88 88 D_lateral AREA=3.125E-016    
M2755 1552 1521 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2754 1520 1527 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2753 88 1524 1526 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2752 1526 1517 1774 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2751 1517 1522 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2750 1525 1522 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2749 1774 1518 1525 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2748 1552 1521 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2747 1520 1527 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2746 1519 1524 1774 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2745 1774 1517 1523 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2744 104 1522 1519 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2743 1517 1522 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2742 1523 1518 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D2741 are shorted:
* D2741 104 104 D_lateral AREA=3.125E-016    $ (-352.5 401.999 -347.5 402)CMOSN2741 104 104 D_lateral AREA=3.125E-016    
M2740 88 1528 1527 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2739 1527 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2738 1527 1528 1529 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2737 1529 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2736 are shorted:
* D2736 88 88 D_lateral AREA=3.125E-016    $ (-416.5 415.5 -416.499 420.5)CMOSN2736 88 88 D_lateral AREA=3.125E-016    
M2735 1538 1530 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2734 1537 1531 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2733 88 1552 1531 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2732 1531 1532 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2731 88 1532 1530 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2730 1530 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2729 1538 1530 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2728 1537 1531 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2727 1531 1552 1534 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2726 1534 1532 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2725 1530 1532 1533 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2724 1533 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2723 are shorted:
* D2723 88 88 D_lateral AREA=3.125E-016    $ (-510 415.5 -509.999 420.5)CMOSN2723 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2722 are shorted:
* D2722 88 88 D_lateral AREA=3.125E-016    $ (-554.5 415.5 -554.499 420.5)CMOSN2722 88 88 D_lateral AREA=3.125E-016    
M2721 1574 1548 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2720 1543 1537 1544 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M2719 88 1538 1543 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M2718 1544 1547 1548 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M2717 1536 1539 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2716 88 1536 1535 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2715 88 1536 1542 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2714 1542 1545 1812 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2713 1541 1549 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2712 1812 1535 1541 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2711 1574 1548 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2710 1548 1537 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M2709 104 1538 1548 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M2708 104 1547 1548 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M2707 1536 1539 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2706 1546 1536 1812 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2705 104 1536 1535 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2704 1812 1545 1540 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2703 1540 1535 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D2702 are shorted:
* D2702 104 104 D_lateral AREA=3.125E-016    $ (-602.501 353.5 -602.5 358.5)CMOSN2702 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2701 are shorted:
* D2701 88 88 D_lateral AREA=3.125E-016    $ (-604 370.5 -603.999 375.5)CMOSN2701 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2700 are shorted:
* D2700 88 88 D_lateral AREA=3.125E-016    $ (-648.5 415.999 -643.5 416)CMOSN2700 88 88 D_lateral AREA=3.125E-016    
M2699 1547 1550 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2698 88 1552 1550 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2697 1545 1549 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2696 1547 1550 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2695 1545 1549 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2694 104 1549 1546 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D2693 are shorted:
* D2693 88 88 D_lateral AREA=3.125E-016    $ (-781 415.5 -780.999 420.5)CMOSN2693 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2692 are shorted:
* D2692 104 104 D_lateral AREA=3.125E-016    $ (-717 401.999 -712 402)CMOSN2692 104 104 D_lateral AREA=3.125E-016    
M2691 1550 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2690 1568 1556 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2689 88 1574 1556 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2687 1553 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2686 1550 1552 1553 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2685 1568 1556 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2684 1556 1574 1551 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
* Pins of element D2682 are shorted:
* D2682 88 88 D_lateral AREA=3.125E-016    $ (-873.5 415.5 -873.499 420.5)CMOSN2682 88 88 D_lateral AREA=3.125E-016    
M2681 1560 1568 1571 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M2680 88 1554 1560 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M2679 1554 1555 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2678 88 1557 1556 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2677 88 1557 1555 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2676 1555 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2675 1564 1558 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2673 104 1554 1565 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M2672 1554 1555 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2671 104 1557 1551 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2670 1555 1557 1559 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2669 1559 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2668 1564 1558 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D2667 are shorted:
* D2667 88 88 D_lateral AREA=3.125E-016    $ (-967.5 370.5 -967.499 375.5)CMOSN2667 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2666 are shorted:
* D2666 104 104 D_lateral AREA=3.125E-016    $ (-966.001 353.5 -966 358.5)CMOSN2666 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2665 are shorted:
* D2665 88 88 D_lateral AREA=3.125E-016    $ (-918 415.5 -917.999 420.5)CMOSN2665 88 88 D_lateral AREA=3.125E-016    
M2664 1596 1565 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2663 1571 1572 1565 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M2662 88 1564 1562 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2661 88 1564 1570 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2660 1570 1561 1851 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2659 1561 1566 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2658 1569 1566 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2657 1851 1562 1569 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2656 1596 1565 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2655 104 1568 1565 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=1.15625p PS=3.5u    
M2654 104 1572 1565 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M2653 1563 1564 1851 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2652 104 1564 1562 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2651 1851 1561 1567 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2650 104 1566 1563 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2649 1561 1566 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2648 1567 1562 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D2647 are shorted:
* D2647 88 88 D_lateral AREA=3.125E-016    $ (-1012 415.999 -1007 416)CMOSN2647 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2646 are shorted:
* D2646 104 104 D_lateral AREA=3.125E-016    $ (-1080.5 401.999 -1075.5 402)CMOSN2646 104 104 D_lateral AREA=3.125E-016    
M2645 1572 1573 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2644 88 1574 1573 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2643 1573 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2642 1572 1573 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2641 1573 1574 1575 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2640 1575 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2639 are shorted:
* D2639 88 88 D_lateral AREA=3.125E-016    $ (-1144.5 415.5 -1144.499 420.5)CMOSN2639 88 88 D_lateral AREA=3.125E-016    
M2638 1578 1576 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2637 88 1596 1576 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2636 1576 1373 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2635 1578 1576 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2634 1576 1596 1577 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2633 1577 1373 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2632 are shorted:
* D2632 88 88 D_lateral AREA=3.125E-016    $ (-1245 415.5 -1244.999 420.5)CMOSN2632 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2631 are shorted:
* D2631 88 88 D_lateral AREA=3.125E-016    $ (-1289.5 415.5 -1289.499 420.5)CMOSN2631 88 88 D_lateral AREA=3.125E-016    
M2630 1583 1578 1584 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M2629 88 1579 1583 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M2628 1584 1588 1589 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M2627 1579 1580 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2626 88 1373 1580 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2625 1580 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2624 1592 1581 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2623 1586 1592 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M2622 1589 1578 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M2621 104 1579 1589 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M2620 104 1588 1589 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M2619 1579 1580 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2618 1580 1373 1582 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2617 1582 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2616 1592 1581 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2615 104 1592 1586 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D2614 are shorted:
* D2614 104 104 D_lateral AREA=3.125E-016    $ (-1337.501 353.5 -1337.5 358.5)CMOSN2614 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2613 are shorted:
* D2613 88 88 D_lateral AREA=3.125E-016    $ (-1339 370.5 -1338.999 375.5)CMOSN2613 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2612 are shorted:
* D2612 88 88 D_lateral AREA=3.125E-016    $ (-1383.5 415.999 -1378.5 416)CMOSN2612 88 88 D_lateral AREA=3.125E-016    
M2611 1619 1589 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2610 1588 1595 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2609 88 1592 1594 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2608 1594 1585 1867 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2607 1585 1590 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2606 1593 1590 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2605 1867 1586 1593 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2604 1619 1589 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2603 1588 1595 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2602 1587 1592 1867 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2601 1867 1585 1591 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2600 104 1590 1587 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2599 1585 1590 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2598 1591 1586 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D2597 are shorted:
* D2597 104 104 D_lateral AREA=3.125E-016    $ (-1452 401.999 -1447 402)CMOSN2597 104 104 D_lateral AREA=3.125E-016    
M2596 88 1596 1595 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2595 1595 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2594 1595 1596 1597 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2593 1597 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2592 are shorted:
* D2592 88 88 D_lateral AREA=3.125E-016    $ (-1516 415.5 -1515.999 420.5)CMOSN2592 88 88 D_lateral AREA=3.125E-016    
M2591 1606 1598 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2590 1605 1599 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2589 88 1619 1599 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2588 1599 1600 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2587 88 1600 1598 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2586 1598 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2585 1606 1598 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2584 1605 1599 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2583 1599 1619 1602 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2582 1602 1600 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2581 1598 1600 1601 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2580 1601 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2579 are shorted:
* D2579 88 88 D_lateral AREA=3.125E-016    $ (-1613 415.5 -1612.999 420.5)CMOSN2579 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2578 are shorted:
* D2578 88 88 D_lateral AREA=3.125E-016    $ (-1657.5 415.5 -1657.499 420.5)CMOSN2578 88 88 D_lateral AREA=3.125E-016    
M2577 1640 1615 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2576 1610 1605 1611 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M2575 88 1606 1610 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M2574 1611 1614 1615 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M2573 1604 1607 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2572 88 1604 1603 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2571 88 1604 1609 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2570 1609 1612 1904 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2569 1904 1603 1616 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2568 1640 1615 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2567 1615 1605 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M2566 104 1606 1615 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M2565 104 1614 1615 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M2564 1604 1607 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2563 1613 1604 1904 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2562 104 1604 1603 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2561 1904 1612 1608 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2560 1608 1603 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D2559 are shorted:
* D2559 104 104 D_lateral AREA=3.125E-016    $ (-1705.501 353.5 -1705.5 358.5)CMOSN2559 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2558 are shorted:
* D2558 88 88 D_lateral AREA=3.125E-016    $ (-1707 370.5 -1706.999 375.5)CMOSN2558 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2557 are shorted:
* D2557 88 88 D_lateral AREA=3.125E-016    $ (-1751.5 415.999 -1746.5 416)CMOSN2557 88 88 D_lateral AREA=3.125E-016    M2556 1614 1617 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2554 1612 1404 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2553 1616 1404 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2552 1614 1617 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2551 1612 1404 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2550 104 1404 1613 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D2549 are shorted:
* D2549 88 88 D_lateral AREA=3.125E-016    $ (-1884 415.5 -1883.999 420.5)CMOSN2549 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2548 are shorted:
* D2548 104 104 D_lateral AREA=3.125E-016    $ (-1820 401.999 -1815 402)CMOSN2548 104 104 D_lateral AREA=3.125E-016    
M2547 1631 1625 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2546 88 1640 1625 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2545 1617 1619 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2544 1617 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2543 1631 1625 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2542 1625 1640 1624 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2541 1617 1619 1618 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2540 1618 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2539 are shorted:
* D2539 88 88 D_lateral AREA=3.125E-016    $ (-1977 415.5 -1976.999 420.5)CMOSN2539 88 88 D_lateral AREA=3.125E-016    
M2538 88 1620 1636 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M2537 1620 1621 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2536 1625 1622 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2535 88 1622 1621 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2534 1621 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2533 1629 1425 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2532 104 1620 1630 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M2530 1620 1621 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2529 1624 1622 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2528 1621 1622 1623 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2527 1623 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2526 1629 1425 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D2525 are shorted:
* D2525 88 88 D_lateral AREA=3.125E-016    $ (-2071 370.5 -2070.999 375.5)CMOSN2525 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2524 are shorted:
* D2524 104 104 D_lateral AREA=3.125E-016    $ (-2069.501 353.5 -2069.5 358.5)CMOSN2524 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2523 are shorted:
* D2523 88 88 D_lateral AREA=3.125E-016    $ (-2021.5 415.5 -2021.499 420.5)CMOSN2523 88 88 D_lateral AREA=3.125E-016    
M2522 1662 1630 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2521 1636 1631 1637 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M2520 1637 1638 1630 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M2519 88 1629 1627 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2518 88 1629 1635 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2517 1635 1626 1933 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2516 1626 1632 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2515 1634 1632 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2514 1933 1627 1634 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2513 1662 1630 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2512 104 1631 1630 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=1.15625p PS=3.5u    
M2511 104 1638 1630 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M2510 1628 1629 1933 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2509 104 1629 1627 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2508 1933 1626 1633 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2507 104 1632 1628 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2506 1626 1632 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2505 1633 1627 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D2504 are shorted:
* D2504 88 88 D_lateral AREA=3.125E-016    $ (-2115.5 415.999 -2110.5 416)CMOSN2504 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2503 are shorted:
* D2503 104 104 D_lateral AREA=3.125E-016    $ (-2184 401.999 -2179 402)CMOSN2503 104 104 D_lateral AREA=3.125E-016    
M2502 1638 1639 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2501 88 1640 1639 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2500 1639 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2499 1638 1639 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2498 1639 1640 1641 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2497 1641 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2496 are shorted:
* D2496 88 88 D_lateral AREA=3.125E-016    $ (-2248 415.5 -2247.999 420.5)CMOSN2496 88 88 D_lateral AREA=3.125E-016    
M2495 1644 1642 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2494 88 1662 1642 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2493 1642 1441 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2492 1644 1642 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2491 1642 1662 1643 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2490 1643 1441 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2489 are shorted:
* D2489 88 88 D_lateral AREA=3.125E-016    $ (-2347.5 415.5 -2347.499 420.5)CMOSN2489 88 88 D_lateral AREA=3.125E-016    
M2488 1649 1644 1650 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M2487 88 1645 1649 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M2486 1650 1654 1655 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M2485 1645 1646 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2484 88 1441 1646 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2483 1646 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2482 1658 1647 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2481 1651 1658 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M2480 1655 1644 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M2479 104 1645 1655 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M2478 104 1654 1655 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M2477 1645 1646 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2476 1646 1441 1648 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2475 1648 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2474 1658 1647 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2473 104 1658 1651 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D2472 are shorted:
* D2472 104 104 D_lateral AREA=3.125E-016    $ (-2440.001 353.5 -2440 358.5)CMOSN2472 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2471 are shorted:
* D2471 88 88 D_lateral AREA=3.125E-016    $ (-2441.5 370.5 -2441.499 375.5)CMOSN2471 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2470 are shorted:
* D2470 88 88 D_lateral AREA=3.125E-016    $ (-2392 415.5 -2391.999 420.5)CMOSN2470 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2469 are shorted:
* D2469 88 88 D_lateral AREA=3.125E-016    $ (-2486 415.999 -2481 416)CMOSN2469 88 88 D_lateral AREA=3.125E-016    
M2468 1683 1655 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2467 1654 1661 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2466 88 1658 1660 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2465 1660 1652 1959 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2464 1652 1656 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2463 1659 1656 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2462 1959 1651 1659 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2461 1683 1655 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2460 1654 1661 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2459 1653 1658 1959 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2458 1959 1652 1657 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2457 104 1656 1653 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2456 1652 1656 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2455 1657 1651 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D2454 are shorted:
* D2454 104 104 D_lateral AREA=3.125E-016    $ (-2554.5 401.999 -2549.5 402)CMOSN2454 104 104 D_lateral AREA=3.125E-016    
M2453 88 1662 1661 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2452 1661 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2451 1661 1662 1663 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2450 1663 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2449 are shorted:
* D2449 88 88 D_lateral AREA=3.125E-016    $ (-2618.5 415.5 -2618.499 420.5)CMOSN2449 88 88 D_lateral AREA=3.125E-016    
M2448 1672 1664 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2447 1671 1665 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2446 88 1683 1665 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2445 1665 1666 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2444 88 1666 1664 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2443 1664 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2442 1672 1664 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2441 1671 1665 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2440 1665 1683 1668 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2439 1668 1666 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2438 1664 1666 1667 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2437 1667 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2436 are shorted:
* D2436 88 88 D_lateral AREA=3.125E-016    $ (-2714.5 415.5 -2714.499 420.5)CMOSN2436 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2435 are shorted:
* D2435 88 88 D_lateral AREA=3.125E-016    $ (-2759 415.5 -2758.999 420.5)CMOSN2435 88 88 D_lateral AREA=3.125E-016    
M2434 1694 1681 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2433 1676 1671 1677 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M2432 88 1672 1676 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M2431 1677 1680 1681 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M2430 1670 1673 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2429 88 1670 1669 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2428 88 1670 1675 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2427 1675 1678 1994 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2426 1994 1669 1682 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2425 1694 1681 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2424 1681 1671 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M2423 104 1672 1681 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M2422 104 1680 1681 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M2421 1670 1673 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2420 1679 1670 1994 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2419 104 1670 1669 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2418 1994 1678 1674 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2417 1674 1669 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D2416 are shorted:
* D2416 104 104 D_lateral AREA=3.125E-016    $ (-2807.001 353.5 -2807 358.5)CMOSN2416 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2415 are shorted:
* D2415 88 88 D_lateral AREA=3.125E-016    $ (-2808.5 370.5 -2808.499 375.5)CMOSN2415 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2414 are shorted:
* D2414 88 88 D_lateral AREA=3.125E-016    $ (-2853 415.999 -2848 416)CMOSN2414 88 88 D_lateral AREA=3.125E-016    
M2413 1680 1684 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2412 1678 1472 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2411 1682 1472 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2410 1680 1684 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2409 1678 1472 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2408 104 1472 1679 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D2407 are shorted:
* D2407 88 88 D_lateral AREA=3.125E-016    $ (-2985.5 415.5 -2985.499 420.5)CMOSN2407 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2406 are shorted:
* D2406 104 104 D_lateral AREA=3.125E-016    $ (-2921.5 401.999 -2916.5 402)CMOSN2406 104 104 D_lateral AREA=3.125E-016    
M2405 88 1683 1684 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2404 1684 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2403 1684 1683 1685 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2402 1685 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2401 88 1349 1686 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2400 88 1349 1691 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2399 1691 1692 2017 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2398 1690 1697 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2397 2017 1686 1690 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2396 1349 1687 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M2395 88 1481 1687 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2394 1687 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2393 1693 1349 2017 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2392 104 1349 1686 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2391 2017 1692 1689 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2390 104 1697 1693 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2389 1689 1686 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M2388 1349 1687 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2387 1687 1481 1688 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2386 1688 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2385 are shorted:
* D2385 88 88 D_lateral AREA=3.125E-016    $ (-3245 369.499 -3240 369.5)CMOSN2385 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2384 are shorted:
* D2384 88 88 D_lateral AREA=3.125E-016    $ (-3268 414 -3267.999 419)CMOSN2384 88 88 D_lateral AREA=3.125E-016    
M2383 1692 1697 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2382 1697 1695 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M2381 88 1694 1695 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2379 1698 1696 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M2378 88 1484 1696 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2377 1696 1701 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2376 1692 1697 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2375 1697 1695 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2374 1695 1694 1700 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2372 1698 1696 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2371 1696 1484 1699 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2370 1699 1701 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2369 are shorted:
* D2369 104 104 D_lateral AREA=3.125E-016    $ (-3313.5 355.499 -3308.5 355.5)CMOSN2369 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2368 are shorted:
* D2368 88 88 D_lateral AREA=3.125E-016    $ (-3373 369 -3372.999 374)CMOSN2368 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2367 are shorted:
* D2367 88 88 D_lateral AREA=3.125E-016    $ (-3352 414 -3351.999 419)CMOSN2367 88 88 D_lateral AREA=3.125E-016    
M2366 88 491 1695 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2365 1701 491 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M2364 104 491 1700 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2363 1701 491 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D2361 are shorted:
* D2361 88 88 D_lateral AREA=3.125E-016    $ (217.5 253 217.501 258)CMOSN2361 88 88 D_lateral AREA=3.125E-016    
M2360 88 1805 1703 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2359 88 1805 1710 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2358 1710 1702 1705 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2357 1702 1717 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2356 1709 1717 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2355 1705 1703 1709 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2354 2020 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2353 2020 1705 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2352 88 1705 2019 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2351 2019 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2350 2023 1718 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2349 88 1721 1718 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2348 1704 1805 1705 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2347 104 1805 1703 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2346 1705 1702 1708 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2345 104 1717 1704 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2344 1702 1717 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2343 1708 1703 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M2342 2020 104 1707 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2341 1707 1705 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2340 2019 1705 1706 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2339 1706 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2338 2023 1718 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D2337 are shorted:
* D2337 88 88 D_lateral AREA=3.125E-016    $ (203 297.499 208 297.5)CMOSN2337 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2336 are shorted:
* D2336 104 104 D_lateral AREA=3.125E-016    $ (134.5 283.499 139.5 283.5)CMOSN2336 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2335 are shorted:
* D2335 88 88 D_lateral AREA=3.125E-016    $ (173 253 173.001 258)CMOSN2335 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2334 are shorted:
* D2334 88 88 D_lateral AREA=3.125E-016    $ (118.5 297 118.501 302)CMOSN2334 88 88 D_lateral AREA=3.125E-016    
M2333 88 1717 1712 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2332 88 1717 1727 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2331 1727 1711 1719 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2330 1711 1728 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2329 1726 1728 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2328 1719 1712 1726 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2327 1718 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2326 88 2023 1715 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2325 88 2023 1725 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2324 1725 1714 2218 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2323 1714 1719 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2322 1724 1719 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2321 2218 1715 1724 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2320 1713 1717 1719 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2319 104 1717 1712 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2318 1719 1711 1723 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2317 104 1728 1713 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2316 1711 1728 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2315 1723 1712 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M2314 1722 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2313 1718 1721 1722 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2312 1716 2023 2218 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2311 104 2023 1715 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2310 2218 1714 1720 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2309 104 1719 1716 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2308 1714 1719 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2307 1720 1715 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D2306 are shorted:
* D2306 88 88 D_lateral AREA=3.125E-016    $ (72.5 297.499 77.5 297.5)CMOSN2306 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2304 are shorted:
* D2304 88 88 D_lateral AREA=3.125E-016    $ (79 253.499 84 253.5)CMOSN2304 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2303 are shorted:
* D2303 104 104 D_lateral AREA=3.125E-016    $ (10.5 239.499 15.5 239.5)CMOSN2303 104 104 D_lateral AREA=3.125E-016    
M2302 88 1729 1728 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2301 1730 2031 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2300 88 104 2031 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2299 2031 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2298 88 1721 1729 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2297 1729 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2296 104 1729 1728 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2295 1730 2031 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2294 2031 104 1732 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2293 1732 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2292 1729 1721 1731 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2291 1731 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2290 are shorted:
* D2290 88 88 D_lateral AREA=3.125E-016    $ (-53.5 253 -53.499 258)CMOSN2290 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2289 are shorted:
* D2289 104 104 D_lateral AREA=3.125E-016    $ (4 283.499 9 283.5)CMOSN2289 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2288 are shorted:
* D2288 88 88 D_lateral AREA=3.125E-016    $ (-53 297 -52.999 302)CMOSN2288 88 88 D_lateral AREA=3.125E-016    
M2287 88 1805 1742 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2286 88 1805 1734 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2285 1734 1739 1741 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2284 88 1761 2032 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2283 2032 1741 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2282 1735 1805 1741 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2281 104 1805 1742 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2279 2032 1761 1733 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2278 1733 1741 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2277 are shorted:
* D2277 88 88 D_lateral AREA=3.125E-016    $ (-160.5 297.499 -155.5 297.5)CMOSN2277 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2276 are shorted:
* D2276 88 88 D_lateral AREA=3.125E-016    $ (-146 253 -145.999 258)CMOSN2276 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2275 are shorted:
* D2275 88 88 D_lateral AREA=3.125E-016    $ (-190.5 253 -190.499 258)CMOSN2275 88 88 D_lateral AREA=3.125E-016    
M2274 1739 1747 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2273 1743 1747 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2272 1741 1742 1743 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2271 88 1741 2036 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2270 2036 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2269 1753 1736 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2268 88 1721 1736 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2267 1736 1761 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2266 1749 1753 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M2265 1740 1739 1741 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=1.84375p PS=4.375u    
M2264 1739 1747 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2263 104 1747 1735 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2262 1740 1742 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M2261 2036 1741 1738 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2260 1738 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2259 1753 1736 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2257 1736 1721 1737 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2256 1737 1761 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2255 104 1753 1749 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D2254 are shorted:
* D2254 104 104 D_lateral AREA=3.125E-016    $ (-229 283.499 -224 283.5)CMOSN2254 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2253 are shorted:
* D2253 88 88 D_lateral AREA=3.125E-016    $ (-291 297.499 -286 297.5)CMOSN2253 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2252 are shorted:
* D2252 88 88 D_lateral AREA=3.125E-016    $ (-245 297 -244.999 302)CMOSN2252 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2251 are shorted:
* D2251 88 88 D_lateral AREA=3.125E-016    $ (-284.5 253.499 -279.5 253.5)CMOSN2251 88 88 D_lateral AREA=3.125E-016    
M2250 88 1759 1760 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2249 2042 2045 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2248 88 1747 1745 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2247 88 1747 1758 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2246 1758 1744 1751 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2245 1744 1760 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2244 1757 1760 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2243 1751 1745 1757 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2242 88 1753 1756 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2241 1756 1748 2257 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2240 1748 1751 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2239 1755 1751 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2238 2257 1749 1755 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2237 104 1759 1760 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2236 2042 2045 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2235 1746 1747 1751 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2234 1745 1747 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2233 1751 1744 1754 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2232 104 1760 1746 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2231 1744 1760 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2230 1754 1745 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M2229 1750 1753 2257 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2228 2257 1748 1752 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2227 104 1751 1750 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2226 1748 1751 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2225 1752 1749 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D2224 are shorted:
* D2224 104 104 D_lateral AREA=3.125E-016    $ (-359.5 283.499 -354.5 283.5)CMOSN2224 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2223 are shorted:
* D2223 104 104 D_lateral AREA=3.125E-016    $ (-353 239.499 -348 239.5)CMOSN2223 104 104 D_lateral AREA=3.125E-016    
M2222 88 1761 2045 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2221 2045 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2220 88 1721 1759 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2219 1759 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2218 2045 1761 1763 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2217 1763 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2216 1759 1721 1762 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2215 1762 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2214 are shorted:
* D2214 88 88 D_lateral AREA=3.125E-016    $ (-417 253 -416.999 258)CMOSN2214 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2213 are shorted:
* D2213 88 88 D_lateral AREA=3.125E-016    $ (-416.5 297 -416.499 302)CMOSN2213 88 88 D_lateral AREA=3.125E-016    
M2212 88 1805 1765 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2211 88 1805 1772 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2210 1772 1764 1767 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2209 1764 1774 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2208 1771 1774 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2207 1767 1765 1771 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2206 88 1793 2047 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2205 2047 1767 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2204 88 1767 2046 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2203 2046 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2202 1766 1805 1767 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2201 104 1805 1765 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2200 1767 1764 1770 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2199 104 1774 1766 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2198 1764 1774 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2197 1770 1765 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M2196 2047 1793 1769 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2195 1769 1767 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2194 2046 1767 1768 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2193 1768 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2192 are shorted:
* D2192 88 88 D_lateral AREA=3.125E-016    $ (-525 297.499 -520 297.5)CMOSN2192 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2190 are shorted:
* D2190 88 88 D_lateral AREA=3.125E-016    $ (-510.5 253 -510.499 258)CMOSN2190 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2189 are shorted:
* D2189 88 88 D_lateral AREA=3.125E-016    $ (-555 253 -554.999 258)CMOSN2189 88 88 D_lateral AREA=3.125E-016    
M2188 2050 1775 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2187 88 1774 1788 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2186 88 1774 1781 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2185 1781 1782 1787 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2184 88 1721 1775 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2183 1775 1793 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2182 88 2050 1773 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2181 88 2050 1780 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2180 1780 1784 2297 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2179 1779 1787 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2178 2297 1773 1779 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2177 2050 1775 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2176 1783 1774 1787 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2175 104 1774 1788 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2174 1787 1782 1778 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2172 1775 1721 1777 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2171 1777 1793 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2170 1785 2050 2297 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2169 104 2050 1773 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2168 2297 1784 1776 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2167 1776 1773 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D2166 are shorted:
* D2166 104 104 D_lateral AREA=3.125E-016    $ (-593.5 283.499 -588.5 283.5)CMOSN2166 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2165 are shorted:
* D2165 88 88 D_lateral AREA=3.125E-016    $ (-655.5 297.499 -650.5 297.5)CMOSN2165 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2164 are shorted:
* D2164 88 88 D_lateral AREA=3.125E-016    $ (-609.5 297 -609.499 302)CMOSN2164 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2163 are shorted:
* D2163 88 88 D_lateral AREA=3.125E-016    $ (-649 253.499 -644 253.5)CMOSN2163 88 88 D_lateral AREA=3.125E-016    
M2162 88 1790 1786 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2161 2056 2060 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2160 88 1793 2060 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2159 1782 1786 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2158 1789 1786 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2157 1787 1788 1789 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2156 88 1721 1790 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2155 1784 1787 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2154 104 1790 1786 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2153 2056 2060 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2152 1782 1786 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2151 104 1786 1783 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2150 104 1788 1778 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=187.5f PS=1.25u    
M2149 1784 1787 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2148 104 1787 1785 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D2147 are shorted:
* D2147 88 88 D_lateral AREA=3.125E-016    $ (-781.5 253 -781.499 258)CMOSN2147 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2146 are shorted:
* D2146 104 104 D_lateral AREA=3.125E-016    $ (-724 283.499 -719 283.5)CMOSN2146 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2145 are shorted:
* D2145 88 88 D_lateral AREA=3.125E-016    $ (-781 297 -780.999 302)CMOSN2145 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2144 are shorted:
* D2144 104 104 D_lateral AREA=3.125E-016    $ (-717.5 239.499 -712.5 239.5)CMOSN2144 104 104 D_lateral AREA=3.125E-016    
M2143 2060 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2142 1790 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2140 88 1822 2063 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2138 1794 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2137 2060 1793 1794 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2136 1792 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2135 1790 1721 1792 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2134 104 1805 1796 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2133 2063 1822 1791 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
* Pins of element D2131 are shorted:
* D2131 88 88 D_lateral AREA=3.125E-016    $ (-888.5 297.499 -883.5 297.5)CMOSN2131 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2130 are shorted:
* D2130 88 88 D_lateral AREA=3.125E-016    $ (-874 253 -873.999 258)CMOSN2130 88 88 D_lateral AREA=3.125E-016    
M2129 1796 1805 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M2128 88 1805 1804 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2127 1804 1795 1798 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2126 1795 1812 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2125 1803 1812 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2124 1798 1796 1803 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2123 88 1798 2063 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2122 88 1798 2062 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2121 2062 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2120 2067 1799 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2119 88 1721 1799 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2117 1797 1805 1798 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2116 1798 1795 1802 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2115 104 1812 1797 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2114 1795 1812 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2113 1802 1796 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M2112 104 1798 1791 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2111 2062 1798 1801 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2110 1801 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2109 2067 1799 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2108 1799 1721 1800 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
* Pins of element D2106 are shorted:
* D2106 104 104 D_lateral AREA=3.125E-016    $ (-957 283.499 -952 283.5)CMOSN2106 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2105 are shorted:
* D2105 88 88 D_lateral AREA=3.125E-016    $ (-918.5 253 -918.499 258)CMOSN2105 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2104 are shorted:
* D2104 88 88 D_lateral AREA=3.125E-016    $ (-973 297 -972.999 302)CMOSN2104 88 88 D_lateral AREA=3.125E-016    
M2103 88 1812 1807 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2102 88 1812 1819 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2101 1819 1806 1813 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2100 1806 1821 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2099 1818 1821 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2098 1813 1807 1818 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2097 88 1822 1799 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2096 88 2067 1810 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2095 88 2067 1817 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2094 1817 1809 2331 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2093 1809 1813 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2092 1816 1813 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2091 2331 1810 1816 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2090 1808 1812 1813 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2089 104 1812 1807 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2088 1813 1806 1815 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2087 104 1821 1808 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2086 1806 1821 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2085 1815 1807 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M2084 104 1822 1800 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2083 1811 2067 2331 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2082 104 2067 1810 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2081 2331 1809 1814 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2080 104 1813 1811 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2079 1809 1813 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2078 1814 1810 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D2077 are shorted:
* D2077 88 88 D_lateral AREA=3.125E-016    $ (-1019 297.499 -1014 297.5)CMOSN2077 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2076 are shorted:
* D2076 104 104 D_lateral AREA=3.125E-016    $ (-1087.5 283.499 -1082.5 283.5)CMOSN2076 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2075 are shorted:
* D2075 88 88 D_lateral AREA=3.125E-016    $ (-1012.5 253.499 -1007.5 253.5)CMOSN2075 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2074 are shorted:
* D2074 104 104 D_lateral AREA=3.125E-016    $ (-1081 239.499 -1076 239.5)CMOSN2074 104 104 D_lateral AREA=3.125E-016    
M2073 88 1820 1821 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2072 1823 2073 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2071 88 1822 2073 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2070 2073 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2069 88 1721 1820 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2068 1820 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2067 104 1820 1821 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2066 1823 2073 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2065 2073 1822 1825 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2064 1825 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2063 1820 1721 1824 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2062 1824 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2061 are shorted:
* D2061 88 88 D_lateral AREA=3.125E-016    $ (-1145 253 -1144.999 258)CMOSN2061 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2060 are shorted:
* D2060 88 88 D_lateral AREA=3.125E-016    $ (-1144.5 297 -1144.499 302)CMOSN2060 88 88 D_lateral AREA=3.125E-016    
M2059 88 1805 1835 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2058 88 1805 1827 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2057 1827 1832 1834 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2056 88 1854 2075 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2055 2075 1834 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2054 1828 1805 1834 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2053 104 1805 1835 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2051 2075 1854 1826 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2050 1826 1834 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D2049 are shorted:
* D2049 88 88 D_lateral AREA=3.125E-016    $ (-1260 297.499 -1255 297.5)CMOSN2049 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2048 are shorted:
* D2048 88 88 D_lateral AREA=3.125E-016    $ (-1245.5 253 -1245.499 258)CMOSN2048 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2047 are shorted:
* D2047 88 88 D_lateral AREA=3.125E-016    $ (-1290 253 -1289.999 258)CMOSN2047 88 88 D_lateral AREA=3.125E-016    
M2046 1832 1851 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2045 1836 1851 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2044 1834 1835 1836 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2043 88 1834 2079 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2042 2079 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2041 1845 1829 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2040 88 1721 1829 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2039 1829 1854 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2038 1841 1845 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M2037 1833 1832 1834 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=1.84375p PS=4.375u    
M2036 1832 1851 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2035 104 1851 1828 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2034 1833 1835 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M2033 2079 1834 1831 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2032 1831 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2031 1845 1829 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2030 104 1851 1838 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2029 1829 1721 1830 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2028 1830 1854 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2027 104 1845 1841 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D2026 are shorted:
* D2026 104 104 D_lateral AREA=3.125E-016    $ (-1328.5 283.499 -1323.5 283.5)CMOSN2026 104 104 D_lateral AREA=3.125E-016    
* Pins of element D2025 are shorted:
* D2025 88 88 D_lateral AREA=3.125E-016    $ (-1390.5 297.499 -1385.5 297.5)CMOSN2025 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2024 are shorted:
* D2024 88 88 D_lateral AREA=3.125E-016    $ (-1344.5 297 -1344.499 302)CMOSN2024 88 88 D_lateral AREA=3.125E-016    
* Pins of element D2023 are shorted:
* D2023 88 88 D_lateral AREA=3.125E-016    $ (-1384 253.499 -1379 253.5)CMOSN2023 88 88 D_lateral AREA=3.125E-016    
M2022 88 1852 1853 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2021 2084 2088 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M2020 88 1851 1838 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M2019 88 1851 1850 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2018 1850 1837 1843 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2017 1837 1853 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2016 1849 1853 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2015 1843 1838 1849 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2014 88 1845 1848 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M2013 1848 1840 2355 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M2012 1840 1843 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2011 1847 1843 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2010 2355 1841 1847 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M2009 104 1852 1853 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2008 2084 2088 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2007 1839 1851 1843 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2006 1843 1837 1846 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2005 104 1853 1839 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2004 1837 1853 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M2003 1846 1838 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M2002 1842 1845 2355 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M2001 2355 1840 1844 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M2000 104 1843 1842 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1999 1840 1843 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1998 1844 1841 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D1997 are shorted:
* D1997 104 104 D_lateral AREA=3.125E-016    $ (-1459 283.499 -1454 283.5)CMOSN1997 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1996 are shorted:
* D1996 104 104 D_lateral AREA=3.125E-016    $ (-1452.5 239.499 -1447.5 239.5)CMOSN1996 104 104 D_lateral AREA=3.125E-016    
M1995 88 1854 2088 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1994 2088 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1993 88 1721 1852 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1992 1852 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1991 2088 1854 1856 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1990 1856 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1989 1852 1721 1855 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1988 1855 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D1987 are shorted:
* D1987 88 88 D_lateral AREA=3.125E-016    $ (-1516.5 253 -1516.499 258)CMOSN1987 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1986 are shorted:
* D1986 88 88 D_lateral AREA=3.125E-016    $ (-1516 297 -1515.999 302)CMOSN1986 88 88 D_lateral AREA=3.125E-016    
M1985 88 1805 1858 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1984 88 1805 1865 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1983 1865 1857 1860 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1982 1857 1867 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1981 1864 1867 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1980 1860 1858 1864 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1979 88 1886 2090 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1978 2090 1860 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1977 88 1860 2089 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1976 2089 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1975 1859 1805 1860 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1974 104 1805 1858 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1973 1860 1857 1863 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1972 104 1867 1859 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1971 1857 1867 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1970 1863 1858 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M1969 2090 1886 1862 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1968 1862 1860 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1967 2089 1860 1861 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1966 1861 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D1965 are shorted:
* D1965 88 88 D_lateral AREA=3.125E-016    $ (-1628 297.499 -1623 297.5)CMOSN1965 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1964 are shorted:
* D1964 88 88 D_lateral AREA=3.125E-016    $ (-1613.5 253 -1613.499 258)CMOSN1964 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1963 are shorted:
* D1963 88 88 D_lateral AREA=3.125E-016    $ (-1658 253 -1657.999 258)CMOSN1963 88 88 D_lateral AREA=3.125E-016    
M1962 2093 1868 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1961 88 1867 1881 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1960 88 1867 1872 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1959 1872 1873 1880 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1958 88 1721 1868 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1957 1868 1886 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1956 88 2093 1866 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1955 88 2093 1871 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1954 1871 1875 2394 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1953 2394 1866 1879 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1952 2093 1868 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1951 1874 1867 1880 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1950 104 1867 1881 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1949 1880 1873 1878 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1948 1868 1721 1870 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1947 1870 1886 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1946 1876 2093 2394 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1945 104 2093 1866 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1944 2394 1875 1869 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1943 1869 1866 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D1942 are shorted:
* D1942 104 104 D_lateral AREA=3.125E-016    $ (-1696.5 283.499 -1691.5 283.5)CMOSN1942 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1941 are shorted:
* D1941 88 88 D_lateral AREA=3.125E-016    $ (-1758.5 297.499 -1753.5 297.5)CMOSN1941 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1940 are shorted:
* D1940 88 88 D_lateral AREA=3.125E-016    $ (-1712.5 297 -1712.499 302)CMOSN1940 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1939 are shorted:
* D1939 88 88 D_lateral AREA=3.125E-016    $ (-1752 253.499 -1747 253.5)CMOSN1939 88 88 D_lateral AREA=3.125E-016    
M1938 88 1883 1877 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1937 2099 2102 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1935 1873 1877 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1934 1882 1877 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1933 1880 1881 1882 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1931 1875 1880 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1930 1879 1880 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1929 104 1883 1877 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1928 2099 2102 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1927 1873 1877 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1926 104 1877 1874 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1925 1878 1881 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M1924 1875 1880 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1923 104 1880 1876 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D1922 are shorted:
* D1922 88 88 D_lateral AREA=3.125E-016    $ (-1884.5 253 -1884.499 258)CMOSN1922 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1921 are shorted:
* D1921 104 104 D_lateral AREA=3.125E-016    $ (-1827 283.499 -1822 283.5)CMOSN1921 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1920 are shorted:
* D1920 88 88 D_lateral AREA=3.125E-016    $ (-1884 297 -1883.999 302)CMOSN1920 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1919 are shorted:
* D1919 104 104 D_lateral AREA=3.125E-016    $ (-1820.5 239.499 -1815.5 239.5)CMOSN1919 104 104 D_lateral AREA=3.125E-016    
M1918 88 1892 1895 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1917 2102 1886 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1916 2102 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1915 1883 1721 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1914 1883 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1911 2102 1886 1885 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1910 1885 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1909 1883 1721 1884 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1908 1884 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D1906 are shorted:
* D1906 88 88 D_lateral AREA=3.125E-016    $ (-1977.5 253 -1977.499 258)CMOSN1906 88 88 D_lateral AREA=3.125E-016    
M1905 88 1805 1888 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1904 88 1805 1897 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1903 1897 1887 1890 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1902 1887 1904 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1901 1896 1904 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1900 1890 1888 1896 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1899 1895 1890 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1898 88 1890 2104 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1897 2104 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1896 2108 1911 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1895 88 1721 1911 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1894 1889 1805 1890 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1893 1888 1805 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1892 1890 1887 1894 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1891 104 1904 1889 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1890 1887 1904 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1889 1894 1888 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M1888 1893 1890 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1887 1893 1892 1895 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1886 2104 1890 1891 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1885 1891 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1884 2108 1911 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1883 1911 1721 1907 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
* Pins of element D1882 are shorted:
* D1882 88 88 D_lateral AREA=3.125E-016    $ (-1992 297.499 -1987 297.5)CMOSN1882 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1881 are shorted:
* D1881 104 104 D_lateral AREA=3.125E-016    $ (-2060.5 283.499 -2055.5 283.5)CMOSN1881 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1880 are shorted:
* D1880 88 88 D_lateral AREA=3.125E-016    $ (-2022 253 -2021.999 258)CMOSN1880 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1879 are shorted:
* D1879 88 88 D_lateral AREA=3.125E-016    $ (-2076.5 297 -2076.499 302)CMOSN1879 88 88 D_lateral AREA=3.125E-016    
M1878 88 1904 1899 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1877 88 1904 1913 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1876 1913 1898 1905 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1875 1898 1915 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1874 1912 1915 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1873 1905 1899 1912 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1872 1911 1892 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1871 88 2108 1902 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1870 88 2108 1910 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1869 1910 1901 2424 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1868 1901 1905 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1867 1909 1905 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1866 2424 1902 1909 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1865 1900 1904 1905 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1864 104 1904 1899 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1863 1905 1898 1908 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1862 104 1915 1900 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1861 1898 1915 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1860 1908 1899 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M1859 1907 1892 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1858 1903 2108 2424 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1857 104 2108 1902 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1856 2424 1901 1906 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1855 104 1905 1903 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1854 1901 1905 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1853 1906 1902 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D1852 are shorted:
* D1852 88 88 D_lateral AREA=3.125E-016    $ (-2122.5 297.499 -2117.5 297.5)CMOSN1852 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1851 are shorted:
* D1851 104 104 D_lateral AREA=3.125E-016    $ (-2191 283.499 -2186 283.5)CMOSN1851 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1850 are shorted:
* D1850 88 88 D_lateral AREA=3.125E-016    $ (-2116 253.499 -2111 253.5)CMOSN1850 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1849 are shorted:
* D1849 104 104 D_lateral AREA=3.125E-016    $ (-2184.5 239.499 -2179.5 239.5)CMOSN1849 104 104 D_lateral AREA=3.125E-016    
M1848 88 1914 1915 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1847 1916 2115 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1846 88 1892 2115 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1845 2115 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1844 88 1721 1914 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1843 1914 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1842 104 1914 1915 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1841 1916 2115 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1840 2115 1892 1918 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1839 1918 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1838 1914 1721 1917 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1837 1917 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D1836 are shorted:
* D1836 88 88 D_lateral AREA=3.125E-016    $ (-2248.5 253 -2248.499 258)CMOSN1836 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1835 are shorted:
* D1835 88 88 D_lateral AREA=3.125E-016    $ (-2248 297 -2247.999 302)CMOSN1835 88 88 D_lateral AREA=3.125E-016    
M1834 88 1805 1928 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1833 88 1805 1920 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1832 1920 1926 1925 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1831 88 1946 2116 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1830 2116 1925 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1829 1921 1805 1925 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1828 104 1805 1928 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1827 2116 1946 1919 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1826 1919 1925 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D1825 are shorted:
* D1825 88 88 D_lateral AREA=3.125E-016    $ (-2362.5 297.499 -2357.5 297.5)CMOSN1825 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1824 are shorted:
* D1824 88 88 D_lateral AREA=3.125E-016    $ (-2348 253 -2347.999 258)CMOSN1824 88 88 D_lateral AREA=3.125E-016    
M1823 1926 1933 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1822 1929 1933 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1821 1925 1928 1929 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1820 88 1925 2120 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1819 2120 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1818 1939 1922 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1817 88 1721 1922 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1816 1922 1946 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1815 1935 1939 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M1814 1925 1926 1927 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1813 104 1933 1921 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1812 1926 1933 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1811 1927 1928 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M1810 2120 1925 1924 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1809 1924 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1808 1939 1922 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1807 1922 1721 1923 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1806 1923 1946 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1805 104 1939 1935 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D1804 are shorted:
* D1804 104 104 D_lateral AREA=3.125E-016    $ (-2431 283.499 -2426 283.5)CMOSN1804 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1803 are shorted:
* D1803 88 88 D_lateral AREA=3.125E-016    $ (-2392.5 253 -2392.499 258)CMOSN1803 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1801 are shorted:
* D1801 88 88 D_lateral AREA=3.125E-016    $ (-2447 297 -2446.999 302)CMOSN1801 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1800 are shorted:
* D1800 88 88 D_lateral AREA=3.125E-016    $ (-2486.5 253.499 -2481.5 253.5)CMOSN1800 88 88 D_lateral AREA=3.125E-016    
M1798 2125 2129 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1797 88 1933 1931 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1796 88 1933 1944 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1795 1944 1930 1937 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1794 1930 1945 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1793 1943 1945 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1792 1937 1931 1943 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1791 88 1939 1942 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1790 1942 1934 2439 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1789 1934 1937 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1788 1941 1937 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1787 2439 1935 1941 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1785 2125 2129 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1784 1932 1933 1937 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1783 104 1933 1931 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1782 1937 1930 1940 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1781 104 1945 1932 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1780 1930 1945 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1779 1940 1931 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M1778 1936 1939 2439 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1777 2439 1934 1938 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1776 104 1937 1936 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1775 1934 1937 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1774 1938 1935 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D1773 are shorted:
* D1773 88 88 D_lateral AREA=3.125E-016    $ (-2493 297.499 -2488 297.5)CMOSN1773 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1772 are shorted:
* D1772 104 104 D_lateral AREA=3.125E-016    $ (-2561.5 283.499 -2556.5 283.5)CMOSN1772 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1771 are shorted:
* D1771 104 104 D_lateral AREA=3.125E-016    $ (-2555 239.499 -2550 239.5)CMOSN1771 104 104 D_lateral AREA=3.125E-016    
M1770 1945 1949 88 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1769 88 1946 2129 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1768 2129 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1767 88 1721 1949 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1766 1949 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1765 1945 1949 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.90625p PS=5.75u    
M1764 2129 1946 1948 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1763 1948 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1762 1949 1721 1947 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1761 1947 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D1760 are shorted:
* D1760 88 88 D_lateral AREA=3.125E-016    $ (-2619 253 -2618.999 258)CMOSN1760 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1759 are shorted:
* D1759 88 88 D_lateral AREA=3.125E-016    $ (-2618.5 297 -2618.499 302)CMOSN1759 88 88 D_lateral AREA=3.125E-016    
M1758 88 1805 1951 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1757 88 1805 1958 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1756 1958 1950 1953 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1755 1950 1959 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1754 1957 1959 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1753 1953 1951 1957 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1752 88 1976 2132 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1751 2132 1953 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1750 88 1953 2131 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1749 2131 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1748 1952 1805 1953 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1747 104 1805 1951 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1746 1953 1950 1956 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1745 104 1959 1952 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1743 1956 1951 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M1742 2132 1976 1955 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1741 1955 1953 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1740 2131 1953 1954 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1739 1954 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D1738 are shorted:
* D1738 88 88 D_lateral AREA=3.125E-016    $ (-2729.5 297.499 -2724.5 297.5)CMOSN1738 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1737 are shorted:
* D1737 88 88 D_lateral AREA=3.125E-016    $ (-2715 253 -2714.999 258)CMOSN1737 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1736 are shorted:
* D1736 88 88 D_lateral AREA=3.125E-016    $ (-2759.5 253 -2759.499 258)CMOSN1736 88 88 D_lateral AREA=3.125E-016    
M1735 2135 1960 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1734 88 1959 1974 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1733 88 1959 1964 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1732 1964 1969 1973 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1731 88 1721 1960 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1730 1960 1976 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1729 88 2135 1971 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1728 88 2135 1963 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1727 1963 1966 2485 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1725 104 1959 1950 104 CMOSN L=500n W=750n AD=2.21875p PD=6.25u AS=1.75p PS=5.5u    
M1724 2135 1960 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1723 1965 1959 1973 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1722 104 1959 1974 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1720 1960 1721 1962 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1719 1962 1976 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1718 1967 2135 2485 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1717 104 2135 1971 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1716 2485 1966 1961 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1715 1961 1971 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D1714 are shorted:
* D1714 104 104 D_lateral AREA=3.125E-016    $ (-2798 283.499 -2793 283.5)CMOSN1714 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1713 are shorted:
* D1713 88 88 D_lateral AREA=3.125E-016    $ (-2860 297.499 -2855 297.5)CMOSN1713 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1712 are shorted:
* D1712 88 88 D_lateral AREA=3.125E-016    $ (-2814 297 -2813.999 302)CMOSN1712 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1711 are shorted:
* D1711 88 88 D_lateral AREA=3.125E-016    $ (-2853.5 253.499 -2848.5 253.5)CMOSN1711 88 88 D_lateral AREA=3.125E-016    
M1710 88 1977 1968 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1709 2141 2145 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1708 1969 1968 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1707 1975 1968 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1706 1973 1974 1975 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1705 1966 1973 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1704 1972 1973 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1703 1972 1971 2485 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1702 104 1977 1968 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1701 2141 2145 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1700 1970 1969 1973 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=1.84375p PS=4.375u    
M1699 1969 1968 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1698 104 1968 1965 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1697 1970 1974 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M1696 1966 1973 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1695 104 1973 1967 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D1694 are shorted:
* D1694 88 88 D_lateral AREA=3.125E-016    $ (-2986 253 -2985.999 258)CMOSN1694 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1693 are shorted:
* D1693 104 104 D_lateral AREA=3.125E-016    $ (-2928.5 283.499 -2923.5 283.5)CMOSN1693 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1692 are shorted:
* D1692 88 88 D_lateral AREA=3.125E-016    $ (-2985.5 297 -2985.499 302)CMOSN1692 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1691 are shorted:
* D1691 104 104 D_lateral AREA=3.125E-016    $ (-2922 239.499 -2917 239.5)CMOSN1691 104 104 D_lateral AREA=3.125E-016    
M1690 88 1976 2145 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1689 2145 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1688 88 1721 1977 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1687 1977 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1686 2145 1976 1979 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1685 1979 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1684 1977 1721 1978 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1683 1978 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D1682 are shorted:
* D1682 88 88 D_lateral AREA=3.125E-016    $ (-3086.5 253 -3086.499 258)CMOSN1682 88 88 D_lateral AREA=3.125E-016    
M1681 88 1805 1981 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1680 88 1805 1988 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1679 1988 1980 1983 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1678 1980 1994 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1677 1987 1994 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1676 1983 1981 1987 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1675 88 2005 2148 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1674 2148 1983 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1673 88 1983 2147 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1672 2147 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1671 2151 1995 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1670 1982 1805 1983 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1669 104 1805 1981 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1668 1983 1980 1986 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1667 104 1994 1982 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1666 1980 1994 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1665 1986 1981 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M1664 2148 2005 1985 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1663 1985 1983 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1662 2147 1983 1984 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1661 1984 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1660 2151 1995 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D1659 are shorted:
* D1659 88 88 D_lateral AREA=3.125E-016    $ (-3101 297.499 -3096 297.5)CMOSN1659 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1658 are shorted:
* D1658 104 104 D_lateral AREA=3.125E-016    $ (-3169.5 283.499 -3164.5 283.5)CMOSN1658 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1657 are shorted:
* D1657 88 88 D_lateral AREA=3.125E-016    $ (-3131 253 -3130.999 258)CMOSN1657 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1656 are shorted:
* D1656 88 88 D_lateral AREA=3.125E-016    $ (-3185.5 297 -3185.499 302)CMOSN1656 88 88 D_lateral AREA=3.125E-016    
M1655 88 1994 1989 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1654 88 1994 2002 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1653 2002 2009 2007 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1652 2009 2004 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1651 2001 2004 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1650 2007 1989 2001 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1649 88 1721 1995 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1648 1995 2005 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1647 88 2151 1992 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1646 88 2151 2000 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1645 2000 1991 2165 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1644 1991 2007 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1643 1999 2007 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1642 2165 1992 1999 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1641 1990 1994 2007 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1640 104 1994 1989 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1639 2007 2009 1998 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1638 104 2004 1990 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1637 1998 1989 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M1636 1995 1721 1997 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1635 1997 2005 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1634 1993 2151 2165 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1633 104 2151 1992 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1632 2165 1991 1996 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1631 104 2007 1993 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1630 1991 2007 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1629 1996 1992 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D1628 are shorted:
* D1628 88 88 D_lateral AREA=3.125E-016    $ (-3231.5 297.499 -3226.5 297.5)CMOSN1628 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1627 are shorted:
* D1627 88 88 D_lateral AREA=3.125E-016    $ (-3225 253.499 -3220 253.5)CMOSN1627 88 88 D_lateral AREA=3.125E-016    
M1625 88 2003 2004 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1624 2006 2158 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1623 88 2005 2158 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1622 2158 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1621 88 1721 2003 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1620 2003 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1619 104 2003 2004 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1618 2006 2158 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1617 2158 2005 2010 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1616 2010 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1615 2009 2004 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1614 2003 1721 2008 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1613 2008 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D1612 are shorted:
* D1612 88 88 D_lateral AREA=3.125E-016    $ (-3357.5 253 -3357.499 258)CMOSN1612 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1611 are shorted:
* D1611 104 104 D_lateral AREA=3.125E-016    $ (-3300 283.499 -3295 283.5)CMOSN1611 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1610 are shorted:
* D1610 88 88 D_lateral AREA=3.125E-016    $ (-3357 297 -3356.999 302)CMOSN1610 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1609 are shorted:
* D1609 104 104 D_lateral AREA=3.125E-016    $ (-3293.5 239.499 -3288.5 239.5)CMOSN1609 104 104 D_lateral AREA=3.125E-016    
M1608 1805 2164 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M1607 88 2017 2164 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1606 2164 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1605 1721 2011 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M1604 2013 491 88 88 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M1603 2011 2166 2013 88 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M1601 1805 2164 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1600 2164 2017 2012 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1599 2012 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1598 1721 2011 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1597 2011 491 104 104 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M1596 104 2166 2011 104 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
* Pins of element D1594 are shorted:
* D1594 88 88 D_lateral AREA=3.125E-016    $ (-3633 251.5 -3632.999 256.5)CMOSN1594 88 88 D_lateral AREA=3.125E-016    
M1593 88 2174 2166 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M1592 88 2177 2174 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1591 2174 2176 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1590 2176 491 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M1589 1717 2014 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M1588 88 2177 2014 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1587 2014 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1586 104 2174 2166 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1585 2174 2177 2016 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1584 2016 2176 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1583 2176 491 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1582 1717 2014 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1581 2014 2177 2015 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1580 2015 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D1579 are shorted:
* D1579 88 88 D_lateral AREA=3.125E-016    $ (-3717 251.5 -3716.999 256.5)CMOSN1579 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1578 are shorted:
* D1578 88 88 D_lateral AREA=3.125E-016    $ (-3746 297 -3745.999 302)CMOSN1578 88 88 D_lateral AREA=3.125E-016    
M1575 88 2074 2181 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1574 88 2074 2022 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1573 2022 2186 2183 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1572 2186 2201 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1571 2021 2201 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1570 2183 2181 2021 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1569 88 2197 2194 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1568 88 2018 2026 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M1567 2018 2019 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1566 88 2020 2025 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1565 104 2018 2024 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M1564 2018 2019 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1563 104 2020 2025 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D1562 are shorted:
* D1562 88 88 D_lateral AREA=3.125E-016    $ (202.5 135.999 207.5 136)CMOSN1562 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1561 are shorted:
* D1561 88 88 D_lateral AREA=3.125E-016    $ (118 135.5 118.001 140.5)CMOSN1561 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1560 are shorted:
* D1560 88 88 D_lateral AREA=3.125E-016    $ (123.5 208 123.501 213)CMOSN1560 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1559 are shorted:
* D1559 104 104 D_lateral AREA=3.125E-016    $ (124.999 191 125 196)CMOSN1559 104 104 D_lateral AREA=3.125E-016    
M1558 88 2201 2188 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1557 88 2201 2029 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1556 2029 2199 2195 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1555 2199 2030 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1554 2028 2030 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1553 2195 2188 2028 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1552 2194 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1551 1761 2024 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1550 2026 2025 2027 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M1549 2027 1730 2024 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M1548 1761 2024 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1547 2024 2025 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M1546 104 1730 2024 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
* Pins of element D1545 are shorted:
* D1545 88 88 D_lateral AREA=3.125E-016    $ (72 135.999 77 136)CMOSN1545 88 88 D_lateral AREA=3.125E-016    
M1544 88 2208 2030 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1543 88 2197 2208 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1542 2208 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D1541 are shorted:
* D1541 88 88 D_lateral AREA=3.125E-016    $ (-53.5 135.5 -53.499 140.5)CMOSN1541 88 88 D_lateral AREA=3.125E-016    
M1540 88 2074 2219 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1539 88 2074 2033 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1538 2033 2214 2039 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1537 2034 2032 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1536 2034 2032 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D1535 are shorted:
* D1535 88 88 D_lateral AREA=3.125E-016    $ (-161 135.999 -156 136)CMOSN1535 88 88 D_lateral AREA=3.125E-016    
M1534 2214 2218 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1533 2040 2218 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1532 2039 2219 2040 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1531 88 2197 2215 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1530 2215 2240 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1529 2037 2034 2038 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M1528 88 2035 2037 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M1527 2038 2042 2041 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M1526 2035 2036 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1525 2041 2034 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M1524 104 2035 2041 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M1523 104 2042 2041 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M1522 2035 2036 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D1520 are shorted:
* D1520 88 88 D_lateral AREA=3.125E-016    $ (-245.5 135.5 -245.499 140.5)CMOSN1520 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1519 are shorted:
* D1519 104 104 D_lateral AREA=3.125E-016    $ (-238.501 191 -238.5 196)CMOSN1519 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1518 are shorted:
* D1518 88 88 D_lateral AREA=3.125E-016    $ (-240 208 -239.999 213)CMOSN1518 88 88 D_lateral AREA=3.125E-016    
M1517 88 2241 2233 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1516 88 2218 2225 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1515 88 2218 2044 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1514 2044 2234 2230 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1513 2234 2233 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1512 2043 2233 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1511 2230 2225 2043 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1510 1793 2041 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1509 1793 2041 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D1508 are shorted:
* D1508 88 88 D_lateral AREA=3.125E-016    $ (-291.5 135.999 -286.5 136)CMOSN1508 88 88 D_lateral AREA=3.125E-016    
M1507 88 2197 2241 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1506 2241 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D1505 are shorted:
* D1505 88 88 D_lateral AREA=3.125E-016    $ (-417 135.5 -416.999 140.5)CMOSN1505 88 88 D_lateral AREA=3.125E-016    
M1504 88 2074 2244 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1503 88 2074 2049 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1502 2049 2249 2246 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1501 2249 2257 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1500 2048 2257 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1499 2246 2244 2048 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1498 2052 2046 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1497 2051 2047 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1496 2052 2046 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1495 2051 2047 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D1494 are shorted:
* D1494 88 88 D_lateral AREA=3.125E-016    $ (-525.5 135.999 -520.5 136)CMOSN1494 88 88 D_lateral AREA=3.125E-016    
M1493 88 2257 2269 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1492 88 2257 2055 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1491 2055 2263 2058 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1490 88 2197 2253 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1489 2253 2274 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1488 1822 2057 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1487 2053 2051 2054 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M1486 88 2052 2053 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M1485 2054 2056 2057 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M1484 1822 2057 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1483 2057 2051 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M1482 104 2052 2057 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M1481 104 2056 2057 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
* Pins of element D1480 are shorted:
* D1480 88 88 D_lateral AREA=3.125E-016    $ (-656 135.999 -651 136)CMOSN1480 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1479 are shorted:
* D1479 88 88 D_lateral AREA=3.125E-016    $ (-610 135.5 -609.999 140.5)CMOSN1479 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1478 are shorted:
* D1478 104 104 D_lateral AREA=3.125E-016    $ (-603.001 191 -603 196)CMOSN1478 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1477 are shorted:
* D1477 88 88 D_lateral AREA=3.125E-016    $ (-604.5 208 -604.499 213)CMOSN1477 88 88 D_lateral AREA=3.125E-016    
M1476 88 2272 2268 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1475 2263 2268 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1474 2059 2268 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1473 2058 2269 2059 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1472 88 2197 2272 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
* Pins of element D1471 are shorted:
* D1471 88 88 D_lateral AREA=3.125E-016    $ (-781.5 135.5 -781.499 140.5)CMOSN1471 88 88 D_lateral AREA=3.125E-016    
M1469 2272 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1468 2069 2063 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1467 2069 2063 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D1466 are shorted:
* D1466 88 88 D_lateral AREA=3.125E-016    $ (-889 135.999 -884 136)CMOSN1466 88 88 D_lateral AREA=3.125E-016    
M1465 2277 2074 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M1464 88 2074 2066 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1463 2066 2283 2279 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1462 2283 2297 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1461 2065 2297 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1460 2279 2277 2065 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1459 88 2197 2280 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1456 88 2061 2064 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M1455 2061 2062 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1453 104 2061 2068 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M1452 2061 2062 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D1451 are shorted:
* D1451 88 88 D_lateral AREA=3.125E-016    $ (-973.5 135.5 -973.499 140.5)CMOSN1451 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1450 are shorted:
* D1450 88 88 D_lateral AREA=3.125E-016    $ (-968 208 -967.999 213)CMOSN1450 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1449 are shorted:
* D1449 104 104 D_lateral AREA=3.125E-016    $ (-966.501 191 -966.5 196)CMOSN1449 104 104 D_lateral AREA=3.125E-016    
M1448 88 2297 2286 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1447 88 2297 2072 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1446 2072 2295 2292 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1445 2295 2294 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1444 2071 2294 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1443 2292 2286 2071 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1442 88 2305 2280 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1441 1854 2068 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1440 2070 2069 2064 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.125p PS=3.75u    
M1439 2070 1823 2068 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M1438 1854 2068 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1437 104 2069 2068 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=1.15625p PS=3.5u    
M1436 104 1823 2068 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
* Pins of element D1435 are shorted:
* D1435 88 88 D_lateral AREA=3.125E-016    $ (-1019.5 135.999 -1014.5 136)CMOSN1435 88 88 D_lateral AREA=3.125E-016    
M1434 88 2304 2294 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1433 88 2197 2304 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1432 2304 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D1431 are shorted:
* D1431 88 88 D_lateral AREA=3.125E-016    $ (-1145 135.5 -1144.999 140.5)CMOSN1431 88 88 D_lateral AREA=3.125E-016    
M1430 88 2074 2082 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1429 88 2074 2076 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1428 2076 2312 2317 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1426 2077 2075 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1425 2077 2075 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D1424 are shorted:
* D1424 88 88 D_lateral AREA=3.125E-016    $ (-1254 135.999 -1249 136)CMOSN1424 88 88 D_lateral AREA=3.125E-016    
M1423 2312 2331 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1422 2083 2331 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1421 2083 2082 2317 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1420 2320 2331 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M1419 88 2197 2314 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1418 2314 2337 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1417 2080 2077 2081 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M1416 88 2078 2080 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M1415 2081 2084 2085 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M1414 2078 2079 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1413 2085 2077 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M1412 104 2078 2085 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M1411 104 2084 2085 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M1410 2078 2079 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D1409 are shorted:
* D1409 88 88 D_lateral AREA=3.125E-016    $ (-1384.5 135.999 -1379.5 136)CMOSN1409 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1408 are shorted:
* D1408 88 88 D_lateral AREA=3.125E-016    $ (-1338.5 135.5 -1338.499 140.5)CMOSN1408 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1407 are shorted:
* D1407 104 104 D_lateral AREA=3.125E-016    $ (-1338.001 191 -1338 196)CMOSN1407 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1406 are shorted:
* D1406 88 88 D_lateral AREA=3.125E-016    $ (-1339.5 208 -1339.499 213)CMOSN1406 88 88 D_lateral AREA=3.125E-016    
M1405 88 2338 2328 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1404 88 2331 2087 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1403 2087 2329 2325 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1402 2329 2328 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1401 2086 2328 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1400 2325 2320 2086 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1399 1886 2085 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1398 1886 2085 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1397 88 2197 2338 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1396 2338 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D1395 are shorted:
* D1395 88 88 D_lateral AREA=3.125E-016    $ (-1510 135.5 -1509.999 140.5)CMOSN1395 88 88 D_lateral AREA=3.125E-016    
M1394 88 2074 2341 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1393 88 2074 2092 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1392 2092 2346 2343 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1391 2346 2355 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1390 2091 2355 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1389 2343 2341 2091 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1388 2095 2089 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1387 2094 2090 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1386 2095 2089 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1385 2094 2090 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D1384 are shorted:
* D1384 88 88 D_lateral AREA=3.125E-016    $ (-1622 135.999 -1617 136)CMOSN1384 88 88 D_lateral AREA=3.125E-016    
M1383 88 2355 2348 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1382 88 2355 2098 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1381 2098 2361 2366 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1380 2366 2348 2101 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1379 88 2197 2351 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1378 2351 2371 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1377 1892 2100 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1376 2096 2094 2097 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M1375 88 2095 2096 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M1374 2097 2099 2100 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M1373 1892 2100 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1372 2100 2094 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M1371 104 2095 2100 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M1370 104 2099 2100 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
* Pins of element D1369 are shorted:
* D1369 88 88 D_lateral AREA=3.125E-016    $ (-1752.5 135.999 -1747.5 136)CMOSN1369 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1368 are shorted:
* D1368 88 88 D_lateral AREA=3.125E-016    $ (-1706.5 135.5 -1706.499 140.5)CMOSN1368 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1367 are shorted:
* D1367 104 104 D_lateral AREA=3.125E-016    $ (-1706.001 191 -1706 196)CMOSN1367 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1366 are shorted:
* D1366 88 88 D_lateral AREA=3.125E-016    $ (-1707.5 208 -1707.499 213)CMOSN1366 88 88 D_lateral AREA=3.125E-016    
M1365 88 2365 2367 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1364 2361 2367 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1363 2101 2367 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1362 88 2197 2365 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
* Pins of element D1361 are shorted:
* D1361 88 88 D_lateral AREA=3.125E-016    $ (-1878 135.5 -1877.999 140.5)CMOSN1361 88 88 D_lateral AREA=3.125E-016    
M1360 2374 2074 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M1359 2365 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1358 2110 1895 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1357 2110 1895 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D1356 are shorted:
* D1356 88 88 D_lateral AREA=3.125E-016    $ (-1986 135.999 -1981 136)CMOSN1356 88 88 D_lateral AREA=3.125E-016    
M1355 88 2074 2106 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1354 2106 2380 2376 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1353 2380 2394 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1352 2105 2394 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1351 2376 2374 2105 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1350 88 2197 2377 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1349 2377 2107 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1348 88 2103 2111 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M1347 2103 2104 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1346 104 2103 2109 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M1344 2103 2104 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D1343 are shorted:
* D1343 88 88 D_lateral AREA=3.125E-016    $ (-2070.5 135.5 -2070.499 140.5)CMOSN1343 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1342 are shorted:
* D1342 88 88 D_lateral AREA=3.125E-016    $ (-2071.5 208 -2071.499 213)CMOSN1342 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1341 are shorted:
* D1341 104 104 D_lateral AREA=3.125E-016    $ (-2070.001 191 -2070 196)CMOSN1341 104 104 D_lateral AREA=3.125E-016    
M1340 88 2394 2383 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1339 88 2394 2114 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1338 2114 2392 2389 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1337 2392 2391 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1336 2113 2391 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1335 2389 2383 2113 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1334 1946 2109 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1333 2111 2110 2112 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M1332 2112 1916 2109 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M1331 1946 2109 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1330 104 2110 2109 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=1.15625p PS=3.5u    
M1329 104 1916 2109 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
* Pins of element D1328 are shorted:
* D1328 88 88 D_lateral AREA=3.125E-016    $ (-2116.5 135.999 -2111.5 136)CMOSN1328 88 88 D_lateral AREA=3.125E-016    
M1327 88 2400 2391 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1326 88 2197 2400 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1325 2400 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D1324 are shorted:
* D1324 88 88 D_lateral AREA=3.125E-016    $ (-2242 135.5 -2241.999 140.5)CMOSN1324 88 88 D_lateral AREA=3.125E-016    
M1323 88 2074 2411 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1322 88 2074 2117 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1321 2117 2407 2123 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1320 2118 2116 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1319 2118 2116 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D1318 are shorted:
* D1318 88 88 D_lateral AREA=3.125E-016    $ (-2356.5 135.999 -2351.5 136)CMOSN1318 88 88 D_lateral AREA=3.125E-016    
M1317 2407 2424 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1316 2124 2424 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1315 2123 2411 2124 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1314 2414 2424 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M1313 88 2197 2408 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1312 2408 2430 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1311 2121 2118 2122 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M1310 88 2119 2121 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M1309 2122 2125 2126 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M1308 2119 2120 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1307 2126 2118 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M1306 104 2119 2126 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M1305 104 2125 2126 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M1304 2119 2120 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D1303 are shorted:
* D1303 88 88 D_lateral AREA=3.125E-016    $ (-2487 135.999 -2482 136)CMOSN1303 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1302 are shorted:
* D1302 88 88 D_lateral AREA=3.125E-016    $ (-2441 135.5 -2440.999 140.5)CMOSN1302 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1301 are shorted:
* D1301 104 104 D_lateral AREA=3.125E-016    $ (-2440.501 191 -2440.5 196)CMOSN1301 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1300 are shorted:
* D1300 88 88 D_lateral AREA=3.125E-016    $ (-2442 208 -2441.999 213)CMOSN1300 88 88 D_lateral AREA=3.125E-016    
M1299 88 2431 2130 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1298 88 2424 2128 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1297 2128 2422 2419 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1296 2422 2130 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1295 2127 2130 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1294 2419 2414 2127 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1293 1976 2126 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1292 1976 2126 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1291 88 2197 2431 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1290 2431 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D1289 are shorted:
* D1289 88 88 D_lateral AREA=3.125E-016    $ (-2612.5 135.5 -2612.499 140.5)CMOSN1289 88 88 D_lateral AREA=3.125E-016    
M1288 88 2074 2434 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1287 88 2074 2134 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1286 2134 2440 2436 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1285 2440 2439 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1284 2133 2439 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1283 2436 2434 2133 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1282 2137 2131 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1281 2136 2132 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1280 2137 2131 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1279 2136 2132 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D1278 are shorted:
* D1278 88 88 D_lateral AREA=3.125E-016    $ (-2723.5 135.999 -2718.5 136)CMOSN1278 88 88 D_lateral AREA=3.125E-016    
M1277 88 2439 2143 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1276 88 2439 2140 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1275 2140 2453 2458 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1273 88 2197 2444 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1272 2444 2463 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1271 2005 2142 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1270 2138 2136 2139 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M1269 88 2137 2138 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M1268 2139 2141 2142 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M1267 2005 2142 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1266 2142 2136 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M1265 104 2137 2142 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M1264 104 2141 2142 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
* Pins of element D1263 are shorted:
* D1263 88 88 D_lateral AREA=3.125E-016    $ (-2854 135.999 -2849 136)CMOSN1263 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1262 are shorted:
* D1262 88 88 D_lateral AREA=3.125E-016    $ (-2808 135.5 -2807.999 140.5)CMOSN1262 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1261 are shorted:
* D1261 104 104 D_lateral AREA=3.125E-016    $ (-2807.501 191 -2807.5 196)CMOSN1261 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1260 are shorted:
* D1260 88 88 D_lateral AREA=3.125E-016    $ (-2809 208 -2808.999 213)CMOSN1260 88 88 D_lateral AREA=3.125E-016    
M1259 88 2457 2459 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1258 2453 2459 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1257 2144 2459 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1256 2144 2143 2458 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1255 88 2197 2457 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
* Pins of element D1254 are shorted:
* D1254 88 88 D_lateral AREA=3.125E-016    $ (-2979.5 135.5 -2979.499 140.5)CMOSN1254 88 88 D_lateral AREA=3.125E-016    
M1253 2457 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1251 88 2074 2465 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1250 88 2074 2150 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1249 2150 2471 2467 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1248 2471 2485 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1247 2149 2485 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1246 2467 2465 2149 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1245 88 2197 2480 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1244 88 2146 2154 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M1243 2146 2147 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1242 2153 2148 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1241 104 2146 2152 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M1240 2146 2147 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1239 2153 2148 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D1238 are shorted:
* D1238 88 88 D_lateral AREA=3.125E-016    $ (-3095 135.999 -3090 136)CMOSN1238 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1237 are shorted:
* D1237 88 88 D_lateral AREA=3.125E-016    $ (-3179.5 135.5 -3179.499 140.5)CMOSN1237 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1236 are shorted:
* D1236 88 88 D_lateral AREA=3.125E-016    $ (-3180.5 208 -3180.499 213)CMOSN1236 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1235 are shorted:
* D1235 104 104 D_lateral AREA=3.125E-016    $ (-3179.001 191 -3179 196)CMOSN1235 104 104 D_lateral AREA=3.125E-016    
M1234 88 2485 2473 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1233 88 2485 2157 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1232 2157 2483 2479 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1231 2483 2491 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1230 2156 2491 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1229 2479 2473 2156 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1228 2480 2495 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1227 2172 2152 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1226 2154 2153 2155 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M1225 2155 2006 2152 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M1224 2172 2152 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1223 2152 2153 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M1222 104 2006 2152 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
* Pins of element D1221 are shorted:
* D1221 88 88 D_lateral AREA=3.125E-016    $ (-3225.5 135.999 -3220.5 136)CMOSN1221 88 88 D_lateral AREA=3.125E-016    
M1220 88 2494 2491 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1219 88 2197 2494 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1218 2494 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D1217 are shorted:
* D1217 88 88 D_lateral AREA=3.125E-016    $ (-3351 135.5 -3350.999 140.5)CMOSN1217 88 88 D_lateral AREA=3.125E-016    
M1216 88 2074 2505 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1215 88 2074 2159 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
* Pins of element D1213 are shorted:
* D1213 88 88 D_lateral AREA=3.125E-016    $ (-3467.5 135.999 -3462.5 136)CMOSN1213 88 88 D_lateral AREA=3.125E-016    
M1212 2506 2501 2159 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1211 2501 2165 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1210 2160 2165 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1209 2506 2505 2160 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1208 88 2197 2502 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1207 2502 2525 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D1206 are shorted:
* D1206 88 88 D_lateral AREA=3.125E-016    $ (-3552 135.5 -3551.999 140.5)CMOSN1206 88 88 D_lateral AREA=3.125E-016    
M1205 88 1805 2162 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1204 88 1805 2171 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1203 2171 2161 2180 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1202 2161 2175 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1201 2170 2175 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1200 2180 2162 2170 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1199 88 2165 2510 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1198 88 2165 2169 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1197 2169 2520 2517 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1196 2520 2519 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1195 2168 2519 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1194 2517 2510 2168 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1193 2163 1805 2180 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1192 104 1805 2162 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1191 2180 2161 2167 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1190 104 2175 2163 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1189 2161 2175 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1188 2167 2162 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D1187 are shorted:
* D1187 88 88 D_lateral AREA=3.125E-016    $ (-3610 206.999 -3605 207)CMOSN1187 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1186 are shorted:
* D1186 104 104 D_lateral AREA=3.125E-016    $ (-3678.5 192.999 -3673.5 193)CMOSN1186 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1185 are shorted:
* D1185 88 88 D_lateral AREA=3.125E-016    $ (-3598 135.999 -3593 136)CMOSN1185 88 88 D_lateral AREA=3.125E-016    
M1184 2175 2173 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M1183 88 2172 2173 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1182 2173 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1181 88 2526 2519 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1180 88 2197 2526 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1179 2526 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1178 2175 2173 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1177 2173 2172 2178 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1176 2178 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D1175 are shorted:
* D1175 88 88 D_lateral AREA=3.125E-016    $ (-3738 206.5 -3737.999 211.5)CMOSN1175 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1174 are shorted:
* D1174 88 88 D_lateral AREA=3.125E-016    $ (-3723.5 135.5 -3723.499 140.5)CMOSN1174 88 88 D_lateral AREA=3.125E-016    
M1173 2197 2533 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M1172 2179 491 88 88 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M1171 2533 2532 2179 88 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M1170 2201 2542 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M1169 88 2540 2542 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1168 2542 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D1167 are shorted:
* D1167 88 88 D_lateral AREA=3.125E-016    $ (-4057 135.5 -4056.999 140.5)CMOSN1167 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1164 are shorted:
* D1164 88 88 D_lateral AREA=3.125E-016    $ (217 91.5 217.001 96.5)CMOSN1164 88 88 D_lateral AREA=3.125E-016    
M1163 88 2549 2204 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M1162 2549 2550 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1161 2559 2551 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1160 2551 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1159 2551 2183 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1158 88 2183 2550 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1157 2550 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1156 2193 2194 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1155 2182 2074 2183 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1154 2183 2186 2187 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1153 2186 2201 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1152 104 2074 2181 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1151 2187 2181 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M1150 104 2201 2182 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1149 104 2549 2558 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M1148 2549 2550 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1147 104 2551 2559 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1146 2551 104 2185 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1145 2185 2183 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1144 2550 2183 2184 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1143 2184 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1142 2193 2194 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D1141 are shorted:
* D1141 104 104 D_lateral AREA=3.125E-016    $ (134 121.999 139 122)CMOSN1141 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1140 are shorted:
* D1140 88 88 D_lateral AREA=3.125E-016    $ (123 46.5 123.001 51.5)CMOSN1140 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1139 are shorted:
* D1139 104 104 D_lateral AREA=3.125E-016    $ (124.499 29.5 124.5 34.5)CMOSN1139 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1138 are shorted:
* D1138 88 88 D_lateral AREA=3.125E-016    $ (172.5 91.5 172.501 96.5)CMOSN1138 88 88 D_lateral AREA=3.125E-016    
M1137 2240 2558 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1136 2204 2559 2205 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M1135 2205 2206 2558 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M1134 88 2193 2191 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1133 88 2193 2203 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1132 2203 2190 2211 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1131 2190 2195 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1130 2202 2195 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1129 2211 2191 2202 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1128 2240 2558 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1127 2558 2559 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M1126 104 2206 2558 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M1125 2189 2201 2195 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1124 2195 2199 2200 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1123 2199 2030 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1122 104 2201 2188 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1121 2200 2188 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M1120 104 2030 2189 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1119 2194 2197 2198 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1118 2198 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1117 2192 2193 2211 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1116 104 2193 2191 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1115 2211 2190 2196 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1114 104 2195 2192 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1113 2190 2195 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1112 2196 2191 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D1111 are shorted:
* D1111 88 88 D_lateral AREA=3.125E-016    $ (78.5 91.999 83.5 92)CMOSN1111 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1110 are shorted:
* D1110 104 104 D_lateral AREA=3.125E-016    $ (10 77.999 15 78)CMOSN1110 104 104 D_lateral AREA=3.125E-016    
M1109 2206 2207 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1108 88 104 2207 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1107 2207 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1106 104 2208 2030 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1105 2206 2207 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1104 2207 104 2210 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1103 2210 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1102 2208 2197 2209 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1101 2209 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D1100 are shorted:
* D1100 88 88 D_lateral AREA=3.125E-016    $ (-54 91.5 -53.999 96.5)CMOSN1100 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1099 are shorted:
* D1099 104 104 D_lateral AREA=3.125E-016    $ (3.5 121.999 8.5 122)CMOSN1099 104 104 D_lateral AREA=3.125E-016    
M1098 2573 2570 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1097 88 2240 2570 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1096 2570 2039 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1095 2213 2074 2039 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1094 104 2074 2219 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1093 2573 2570 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1092 2570 2240 2212 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1091 2212 2039 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D1090 are shorted:
* D1090 88 88 D_lateral AREA=3.125E-016    $ (-146.5 91.5 -146.499 96.5)CMOSN1090 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1089 are shorted:
* D1089 88 88 D_lateral AREA=3.125E-016    $ (-191 91.5 -190.999 96.5)CMOSN1089 88 88 D_lateral AREA=3.125E-016    
M1088 2221 2573 2222 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M1087 88 2574 2221 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M1086 2222 2229 2223 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M1085 2574 2575 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1084 88 2039 2575 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1083 2575 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1082 2232 2215 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1081 2224 2232 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M1080 2039 2214 2220 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1079 2214 2218 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1078 2220 2219 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M1077 104 2218 2213 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1076 2223 2573 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M1075 104 2574 2223 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M1074 104 2229 2223 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M1073 2574 2575 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1072 2575 2039 2217 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1071 2217 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1070 2232 2215 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1068 2215 2197 2216 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1067 2216 2240 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1066 104 2232 2224 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D1065 are shorted:
* D1065 104 104 D_lateral AREA=3.125E-016    $ (-229.5 121.999 -224.5 122)CMOSN1065 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1064 are shorted:
* D1064 104 104 D_lateral AREA=3.125E-016    $ (-239.001 29.5 -239 34.5)CMOSN1064 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1063 are shorted:
* D1063 88 88 D_lateral AREA=3.125E-016    $ (-240.5 46.5 -240.499 51.5)CMOSN1063 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1062 are shorted:
* D1062 88 88 D_lateral AREA=3.125E-016    $ (-285 91.999 -280 92)CMOSN1062 88 88 D_lateral AREA=3.125E-016    
M1061 2274 2223 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1060 2229 2239 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1059 88 2232 2237 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1058 2237 2227 2238 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1057 2227 2230 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1056 2236 2230 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1055 2238 2224 2236 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1054 104 2241 2233 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1053 2274 2223 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1052 2229 2239 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1051 2226 2218 2230 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1050 2230 2234 2235 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1049 2234 2233 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1048 2225 2218 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1047 2235 2225 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M1046 104 2233 2226 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1045 2228 2232 2238 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1044 2238 2227 2231 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1043 104 2230 2228 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1042 2227 2230 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1041 2231 2224 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D1040 are shorted:
* D1040 104 104 D_lateral AREA=3.125E-016    $ (-360 121.999 -355 122)CMOSN1040 104 104 D_lateral AREA=3.125E-016    
* Pins of element D1039 are shorted:
* D1039 104 104 D_lateral AREA=3.125E-016    $ (-353.5 77.999 -348.5 78)CMOSN1039 104 104 D_lateral AREA=3.125E-016    
M1038 88 2240 2239 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1037 2239 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1036 2239 2240 2243 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1035 2243 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1034 2241 2197 2242 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1033 2242 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D1032 are shorted:
* D1032 88 88 D_lateral AREA=3.125E-016    $ (-417.5 91.5 -417.499 96.5)CMOSN1032 88 88 D_lateral AREA=3.125E-016    
M1031 2603 2597 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1030 2602 2598 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1029 88 2274 2598 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1028 2598 2246 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1027 88 2246 2597 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1026 2597 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1025 2245 2074 2246 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M1024 2246 2249 2250 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M1023 2249 2257 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M1022 104 2074 2244 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1021 2250 2244 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M1020 104 2257 2245 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1019 2603 2597 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1018 2602 2598 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M1017 2598 2274 2248 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1016 2248 2246 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1015 2597 2246 2247 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1014 2247 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D1012 are shorted:
* D1012 88 88 D_lateral AREA=3.125E-016    $ (-511 91.5 -510.999 96.5)CMOSN1012 88 88 D_lateral AREA=3.125E-016    
* Pins of element D1011 are shorted:
* D1011 88 88 D_lateral AREA=3.125E-016    $ (-555.5 91.5 -555.499 96.5)CMOSN1011 88 88 D_lateral AREA=3.125E-016    
M1010 2305 2267 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1009 2260 2602 2261 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M1008 88 2603 2260 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M1007 2261 2266 2267 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M1006 2252 2253 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M1005 88 2252 2251 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M1004 88 2252 2259 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M1003 2259 2264 2270 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M1001 2270 2251 2258 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M1000 2305 2267 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M999 2267 2602 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M998 104 2603 2267 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M997 104 2266 2267 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M996 2252 2253 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M995 2262 2257 2058 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M994 2058 2263 2256 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M993 104 2257 2269 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M991 2253 2197 2255 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M990 2255 2274 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M989 2265 2252 2270 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M988 104 2252 2251 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M987 2270 2264 2254 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M986 2254 2251 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D985 are shorted:
* D985 104 104 D_lateral AREA=3.125E-016    $ (-594 121.999 -589 122)CMOSN985 104 104 D_lateral AREA=3.125E-016    
* Pins of element D984 are shorted:
* D984 104 104 D_lateral AREA=3.125E-016    $ (-603.501 29.5 -603.5 34.5)CMOSN984 104 104 D_lateral AREA=3.125E-016    
* Pins of element D983 are shorted:
* D983 88 88 D_lateral AREA=3.125E-016    $ (-605 46.5 -604.999 51.5)CMOSN983 88 88 D_lateral AREA=3.125E-016    
* Pins of element D982 are shorted:
* D982 88 88 D_lateral AREA=3.125E-016    $ (-649.5 91.999 -644.5 92)CMOSN982 88 88 D_lateral AREA=3.125E-016    
M981 2266 2271 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M980 88 2274 2271 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M979 2264 2058 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M978 88 2058 2258 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M977 104 2272 2268 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M976 2266 2271 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M975 2263 2268 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M974 104 2269 2256 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=187.5f PS=1.25u    
M973 104 2268 2262 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M972 2264 2058 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M971 104 2058 2265 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D970 are shorted:
* D970 88 88 D_lateral AREA=3.125E-016    $ (-782 91.5 -781.999 96.5)CMOSN970 88 88 D_lateral AREA=3.125E-016    
* Pins of element D969 are shorted:
* D969 104 104 D_lateral AREA=3.125E-016    $ (-724.5 121.999 -719.5 122)CMOSN969 104 104 D_lateral AREA=3.125E-016    
* Pins of element D968 are shorted:
* D968 104 104 D_lateral AREA=3.125E-016    $ (-718 77.999 -713 78)CMOSN968 104 104 D_lateral AREA=3.125E-016    
M967 2300 2622 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M966 88 2305 2622 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M964 2271 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M963 104 2074 2277 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M962 2300 2622 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M961 2622 2305 2276 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M959 2271 2274 2275 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M958 2275 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M957 2272 2197 2273 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M956 2273 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D955 are shorted:
* D955 88 88 D_lateral AREA=3.125E-016    $ (-874.5 91.5 -874.499 96.5)CMOSN955 88 88 D_lateral AREA=3.125E-016    
M953 88 2620 2285 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M952 2620 2621 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M951 88 2279 2622 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M950 88 2279 2621 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M949 2621 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M948 2291 2280 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M947 2278 2074 2279 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M946 2279 2283 2284 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M945 2283 2297 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M944 2284 2277 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M943 104 2297 2278 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M941 104 2620 2630 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M940 2620 2621 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M939 104 2279 2276 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M938 2621 2279 2282 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M937 2282 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M936 2291 2280 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M935 2280 2197 2281 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
* Pins of element D933 are shorted:
* D933 104 104 D_lateral AREA=3.125E-016    $ (-957.5 121.999 -952.5 122)CMOSN933 104 104 D_lateral AREA=3.125E-016    
* Pins of element D932 are shorted:
* D932 88 88 D_lateral AREA=3.125E-016    $ (-968.5 46.5 -968.499 51.5)CMOSN932 88 88 D_lateral AREA=3.125E-016    
* Pins of element D931 are shorted:
* D931 104 104 D_lateral AREA=3.125E-016    $ (-967.001 29.5 -967 34.5)CMOSN931 104 104 D_lateral AREA=3.125E-016    
* Pins of element D930 are shorted:
* D930 88 88 D_lateral AREA=3.125E-016    $ (-919 91.5 -918.999 96.5)CMOSN930 88 88 D_lateral AREA=3.125E-016    
M929 2337 2630 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M928 2301 2300 2285 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.125p PS=3.75u    
M927 2301 2302 2630 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M926 88 2291 2289 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M925 88 2291 2299 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M924 2299 2288 2308 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M923 2288 2292 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M922 2298 2292 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M921 2308 2289 2298 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M920 2337 2630 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M919 104 2300 2630 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=1.15625p PS=3.5u    
M918 104 2302 2630 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M917 2287 2297 2292 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M916 2292 2295 2296 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M915 2295 2294 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M914 104 2297 2286 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M913 2296 2286 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M912 104 2294 2287 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M911 104 2305 2281 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M910 2290 2291 2308 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M909 104 2291 2289 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M908 2308 2288 2293 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M907 104 2292 2290 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M906 2288 2292 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M905 2293 2289 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D904 are shorted:
* D904 104 104 D_lateral AREA=3.125E-016    $ (-1088 121.999 -1083 122)CMOSN904 104 104 D_lateral AREA=3.125E-016    
* Pins of element D903 are shorted:
* D903 88 88 D_lateral AREA=3.125E-016    $ (-1013 91.999 -1008 92)CMOSN903 88 88 D_lateral AREA=3.125E-016    
* Pins of element D902 are shorted:
* D902 104 104 D_lateral AREA=3.125E-016    $ (-1081.5 77.999 -1076.5 78)CMOSN902 104 104 D_lateral AREA=3.125E-016    
M901 2302 2303 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M900 88 2305 2303 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M899 2303 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M898 104 2304 2294 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M897 2302 2303 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M896 2303 2305 2307 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M895 2307 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M894 2304 2197 2306 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M893 2306 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D892 are shorted:
* D892 88 88 D_lateral AREA=3.125E-016    $ (-1145.5 91.5 -1145.499 96.5)CMOSN892 88 88 D_lateral AREA=3.125E-016    
M891 2640 2639 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M890 88 2337 2639 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M889 2639 2317 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M887 2311 2074 2317 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M886 2317 2312 2310 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M885 104 2074 2082 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M884 2310 2082 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M883 2640 2639 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M882 2639 2337 2309 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M881 2309 2317 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D880 are shorted:
* D880 88 88 D_lateral AREA=3.125E-016    $ (-1239.5 91.5 -1239.499 96.5)CMOSN880 88 88 D_lateral AREA=3.125E-016    
* Pins of element D879 are shorted:
* D879 88 88 D_lateral AREA=3.125E-016    $ (-1284 91.5 -1283.999 96.5)CMOSN879 88 88 D_lateral AREA=3.125E-016    
M878 2318 2640 2319 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M877 88 2313 2318 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M876 2319 2324 2645 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M875 2313 2643 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M874 2643 2317 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M873 2643 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M872 2327 2314 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M871 2332 2327 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M870 2312 2331 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M869 104 2331 2311 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M868 2645 2640 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M867 104 2313 2645 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M866 104 2324 2645 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M865 2313 2643 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M864 2643 2317 2316 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M863 2316 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M862 2327 2314 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M861 104 2331 2320 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M860 2314 2197 2315 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M859 2315 2337 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M858 104 2327 2332 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D857 are shorted:
* D857 104 104 D_lateral AREA=3.125E-016    $ (-1322.5 121.999 -1317.5 122)CMOSN857 104 104 D_lateral AREA=3.125E-016    
* Pins of element D856 are shorted:
* D856 104 104 D_lateral AREA=3.125E-016    $ (-1332.001 29.5 -1332 34.5)CMOSN856 104 104 D_lateral AREA=3.125E-016    
* Pins of element D855 are shorted:
* D855 88 88 D_lateral AREA=3.125E-016    $ (-1333.5 46.5 -1333.499 51.5)CMOSN855 88 88 D_lateral AREA=3.125E-016    
* Pins of element D854 are shorted:
* D854 88 88 D_lateral AREA=3.125E-016    $ (-1378 91.999 -1373 92)CMOSN854 88 88 D_lateral AREA=3.125E-016    
M853 2371 2645 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M852 2324 2336 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M851 88 2327 2334 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M850 2334 2322 2335 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M849 2322 2325 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M848 2333 2325 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M847 2335 2332 2333 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M846 104 2338 2328 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M845 2371 2645 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M844 2324 2336 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M843 2321 2331 2325 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M842 2325 2329 2330 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M841 2329 2328 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M840 2330 2320 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M839 104 2328 2321 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M838 2323 2327 2335 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M837 2335 2322 2326 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M836 104 2325 2323 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M835 2322 2325 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M834 2326 2332 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D833 are shorted:
* D833 104 104 D_lateral AREA=3.125E-016    $ (-1453 121.999 -1448 122)CMOSN833 104 104 D_lateral AREA=3.125E-016    
* Pins of element D832 are shorted:
* D832 104 104 D_lateral AREA=3.125E-016    $ (-1446.5 77.999 -1441.5 78)CMOSN832 104 104 D_lateral AREA=3.125E-016    
M831 88 2337 2336 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M830 2336 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M829 2336 2337 2340 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M828 2340 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M827 2338 2197 2339 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M826 2339 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D825 are shorted:
* D825 88 88 D_lateral AREA=3.125E-016    $ (-1510.5 91.5 -1510.499 96.5)CMOSN825 88 88 D_lateral AREA=3.125E-016    
M824 2650 2646 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M823 2649 2647 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M822 88 2371 2647 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M821 2647 2343 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M820 88 2343 2646 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M819 2646 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M818 2342 2074 2343 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M817 2343 2346 2347 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M816 2346 2355 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M815 104 2074 2341 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M814 2347 2341 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M813 104 2355 2342 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M812 2650 2646 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M811 2649 2647 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M810 2647 2371 2345 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M809 2345 2343 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M808 2646 2343 2344 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M807 2344 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D806 are shorted:
* D806 104 104 D_lateral AREA=3.125E-016    $ (-1690.5 121.999 -1685.5 122)CMOSN806 104 104 D_lateral AREA=3.125E-016    
* Pins of element D805 are shorted:
* D805 88 88 D_lateral AREA=3.125E-016    $ (-1607.5 91.5 -1607.499 96.5)CMOSN805 88 88 D_lateral AREA=3.125E-016    
* Pins of element D804 are shorted:
* D804 88 88 D_lateral AREA=3.125E-016    $ (-1652 91.5 -1651.999 96.5)CMOSN804 88 88 D_lateral AREA=3.125E-016    
M803 2107 2648 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M802 2358 2649 2359 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M801 88 2650 2358 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M800 2359 2364 2648 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M799 2350 2351 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M798 88 2350 2349 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M797 88 2350 2357 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M796 2357 2362 2368 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M795 2356 2366 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M794 2368 2349 2356 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M793 2107 2648 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M792 2648 2649 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M791 104 2650 2648 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M790 104 2364 2648 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M789 2350 2351 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M788 2360 2355 2366 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M787 2366 2361 2354 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M786 104 2355 2348 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M785 2354 2348 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M784 2351 2197 2353 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M783 2353 2371 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M782 2363 2350 2368 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M781 104 2350 2349 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M780 2368 2362 2352 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M778 2352 2349 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D777 are shorted:
* D777 104 104 D_lateral AREA=3.125E-016    $ (-1700.001 29.5 -1700 34.5)CMOSN777 104 104 D_lateral AREA=3.125E-016    
* Pins of element D776 are shorted:
* D776 88 88 D_lateral AREA=3.125E-016    $ (-1701.5 46.5 -1701.499 51.5)CMOSN776 88 88 D_lateral AREA=3.125E-016    
* Pins of element D775 are shorted:
* D775 88 88 D_lateral AREA=3.125E-016    $ (-1746 91.999 -1741 92)CMOSN775 88 88 D_lateral AREA=3.125E-016    
M774 2364 2369 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M773 88 2371 2369 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M772 2362 2366 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M771 104 2365 2367 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M770 2364 2369 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M768 2361 2367 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M767 104 2367 2360 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M765 2362 2366 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M764 2363 2366 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
* Pins of element D763 are shorted:
* D763 88 88 D_lateral AREA=3.125E-016    $ (-1878.5 91.5 -1878.499 96.5)CMOSN763 88 88 D_lateral AREA=3.125E-016    
* Pins of element D762 are shorted:
* D762 104 104 D_lateral AREA=3.125E-016    $ (-1821 121.999 -1816 122)CMOSN762 104 104 D_lateral AREA=3.125E-016    
* Pins of element D761 are shorted:
* D761 104 104 D_lateral AREA=3.125E-016    $ (-1814.5 77.999 -1809.5 78)CMOSN761 104 104 D_lateral AREA=3.125E-016    
M760 2655 2651 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M759 88 2107 2651 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M758 2651 2376 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M757 2369 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M756 104 2074 2374 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M755 2655 2651 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M754 2651 2107 2373 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M753 2373 2376 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M752 2372 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M751 2372 2371 2369 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M750 2370 2197 2365 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M749 2370 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D748 are shorted:
* D748 88 88 D_lateral AREA=3.125E-016    $ (-1971.5 91.5 -1971.499 96.5)CMOSN748 88 88 D_lateral AREA=3.125E-016    
M747 2382 2655 2397 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M746 88 2652 2382 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M745 2652 2653 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M744 88 2376 2653 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M743 2653 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M742 2388 2377 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M741 2375 2074 2376 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M740 2376 2380 2381 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M739 2380 2394 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M738 2381 2374 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M737 104 2394 2375 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M736 2654 2655 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M735 104 2652 2654 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M734 2652 2653 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M733 2653 2376 2379 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M732 2379 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M731 2388 2377 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M730 2377 2197 2378 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M729 2378 2107 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D728 are shorted:
* D728 104 104 D_lateral AREA=3.125E-016    $ (-2054.5 121.999 -2049.5 122)CMOSN728 104 104 D_lateral AREA=3.125E-016    
* Pins of element D727 are shorted:
* D727 88 88 D_lateral AREA=3.125E-016    $ (-2065.5 46.5 -2065.499 51.5)CMOSN727 88 88 D_lateral AREA=3.125E-016    
* Pins of element D726 are shorted:
* D726 104 104 D_lateral AREA=3.125E-016    $ (-2064.001 29.5 -2064 34.5)CMOSN726 104 104 D_lateral AREA=3.125E-016    
* Pins of element D725 are shorted:
* D725 88 88 D_lateral AREA=3.125E-016    $ (-2016 91.5 -2015.999 96.5)CMOSN725 88 88 D_lateral AREA=3.125E-016    
M724 2430 2654 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M723 2397 2398 2654 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M722 88 2388 2386 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M721 88 2388 2396 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M720 2396 2385 2403 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M719 2385 2389 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M718 2395 2389 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M717 2403 2386 2395 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M716 2430 2654 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M715 104 2398 2654 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M714 2384 2394 2389 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M713 2389 2392 2393 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M712 2392 2391 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M711 104 2394 2383 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M710 2393 2383 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M709 104 2391 2384 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M708 2387 2388 2403 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M707 104 2388 2386 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M706 2403 2385 2390 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M705 104 2389 2387 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M704 2385 2389 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M703 2390 2386 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D702 are shorted:
* D702 104 104 D_lateral AREA=3.125E-016    $ (-2185 121.999 -2180 122)CMOSN702 104 104 D_lateral AREA=3.125E-016    
* Pins of element D701 are shorted:
* D701 88 88 D_lateral AREA=3.125E-016    $ (-2110 91.999 -2105 92)CMOSN701 88 88 D_lateral AREA=3.125E-016    
* Pins of element D700 are shorted:
* D700 104 104 D_lateral AREA=3.125E-016    $ (-2178.5 77.999 -2173.5 78)CMOSN700 104 104 D_lateral AREA=3.125E-016    
M699 2398 2399 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M698 88 2107 2399 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M697 2399 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M696 104 2400 2391 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M695 2398 2399 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M694 2399 2107 2402 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M693 2402 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M692 2400 2197 2401 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M691 2401 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D690 are shorted:
* D690 88 88 D_lateral AREA=3.125E-016    $ (-2242.5 91.5 -2242.499 96.5)CMOSN690 88 88 D_lateral AREA=3.125E-016    
M689 2657 2656 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M688 88 2430 2656 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M687 2656 2123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M686 2406 2074 2123 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M685 2123 2407 2405 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M684 104 2074 2411 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M682 2657 2656 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M681 2656 2430 2404 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M680 2404 2123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D679 are shorted:
* D679 88 88 D_lateral AREA=3.125E-016    $ (-2342 91.5 -2341.999 96.5)CMOSN679 88 88 D_lateral AREA=3.125E-016    
* Pins of element D678 are shorted:
* D678 88 88 D_lateral AREA=3.125E-016    $ (-2386.5 91.5 -2386.499 96.5)CMOSN678 88 88 D_lateral AREA=3.125E-016    
M677 2412 2657 2413 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M676 88 2658 2412 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M675 2413 2418 2660 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M674 2658 2659 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M673 88 2123 2659 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M672 2659 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M671 2421 2408 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M670 2425 2421 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M669 2407 2424 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M668 104 2411 2405 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=187.5f PS=1.25u    
M667 104 2424 2406 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M666 2660 2657 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M665 104 2658 2660 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M664 104 2418 2660 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M663 2658 2659 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M662 2659 2123 2410 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M661 2410 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M660 2421 2408 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M659 104 2424 2414 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M658 2408 2197 2409 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M657 2409 2430 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M656 104 2421 2425 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D655 are shorted:
* D655 104 104 D_lateral AREA=3.125E-016    $ (-2425 121.999 -2420 122)CMOSN655 104 104 D_lateral AREA=3.125E-016    
* Pins of element D654 are shorted:
* D654 104 104 D_lateral AREA=3.125E-016    $ (-2434.501 29.5 -2434.5 34.5)CMOSN654 104 104 D_lateral AREA=3.125E-016    
* Pins of element D653 are shorted:
* D653 88 88 D_lateral AREA=3.125E-016    $ (-2436 46.5 -2435.999 51.5)CMOSN653 88 88 D_lateral AREA=3.125E-016    
* Pins of element D652 are shorted:
* D652 88 88 D_lateral AREA=3.125E-016    $ (-2480.5 91.999 -2475.5 92)CMOSN652 88 88 D_lateral AREA=3.125E-016    
M651 2463 2660 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M650 2418 2429 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M649 88 2421 2427 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M648 2427 2416 2428 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M647 2416 2419 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M646 2426 2419 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M645 2428 2425 2426 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M644 104 2431 2130 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M643 2463 2660 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M642 2418 2429 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M641 2415 2424 2419 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M640 2419 2422 2423 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M639 2422 2130 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M638 2423 2414 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M637 104 2130 2415 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M636 2417 2421 2428 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M635 2428 2416 2420 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M634 104 2419 2417 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M633 2416 2419 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M632 2420 2425 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D631 are shorted:
* D631 104 104 D_lateral AREA=3.125E-016    $ (-2555.5 121.999 -2550.5 122)CMOSN631 104 104 D_lateral AREA=3.125E-016    
* Pins of element D630 are shorted:
* D630 104 104 D_lateral AREA=3.125E-016    $ (-2549 77.999 -2544 78)CMOSN630 104 104 D_lateral AREA=3.125E-016    
M629 88 2430 2429 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M628 2429 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M627 2429 2430 2433 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M626 2433 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M625 2431 2197 2432 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M624 2432 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D623 are shorted:
* D623 88 88 D_lateral AREA=3.125E-016    $ (-2613 91.5 -2612.999 96.5)CMOSN623 88 88 D_lateral AREA=3.125E-016    
M622 2665 2661 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M621 2664 2662 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M620 88 2463 2662 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M619 2662 2436 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M618 88 2436 2661 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M617 2661 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M616 2435 2074 2436 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M615 2436 2440 2441 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M614 2440 2439 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M613 104 2074 2434 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M612 2441 2434 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M611 104 2439 2435 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M610 2665 2661 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M609 2664 2662 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M608 2662 2463 2438 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M607 2438 2436 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M606 2661 2436 2437 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M605 2437 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D603 are shorted:
* D603 88 88 D_lateral AREA=3.125E-016    $ (-2709 91.5 -2708.999 96.5)CMOSN603 88 88 D_lateral AREA=3.125E-016    
* Pins of element D602 are shorted:
* D602 88 88 D_lateral AREA=3.125E-016    $ (-2753.5 91.5 -2753.499 96.5)CMOSN602 88 88 D_lateral AREA=3.125E-016    
M601 2495 2663 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M600 2450 2664 2451 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M599 88 2665 2450 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M598 2451 2456 2663 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M597 2443 2444 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M596 88 2443 2442 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M595 88 2443 2449 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M594 2449 2454 2460 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M593 2448 2458 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M592 2460 2442 2448 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M591 2495 2663 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M590 2663 2664 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M589 104 2665 2663 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M588 104 2456 2663 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M587 2443 2444 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M586 2452 2439 2458 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M585 2458 2453 2447 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M584 104 2439 2143 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M583 2447 2143 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M582 2444 2197 2446 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M581 2446 2463 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M580 2455 2443 2460 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M579 104 2443 2442 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M578 2460 2454 2445 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M576 2445 2442 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D575 are shorted:
* D575 104 104 D_lateral AREA=3.125E-016    $ (-2792 121.999 -2787 122)CMOSN575 104 104 D_lateral AREA=3.125E-016    
* Pins of element D574 are shorted:
* D574 104 104 D_lateral AREA=3.125E-016    $ (-2801.501 29.5 -2801.5 34.5)CMOSN574 104 104 D_lateral AREA=3.125E-016    
* Pins of element D573 are shorted:
* D573 88 88 D_lateral AREA=3.125E-016    $ (-2803 46.5 -2802.999 51.5)CMOSN573 88 88 D_lateral AREA=3.125E-016    
* Pins of element D572 are shorted:
* D572 88 88 D_lateral AREA=3.125E-016    $ (-2847.5 91.999 -2842.5 92)CMOSN572 88 88 D_lateral AREA=3.125E-016    
M571 2456 2461 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M570 88 2463 2461 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M569 2454 2458 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M568 104 2457 2459 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M567 2456 2461 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M565 2453 2459 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M564 104 2459 2452 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M562 2454 2458 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M561 2455 2458 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
* Pins of element D560 are shorted:
* D560 88 88 D_lateral AREA=3.125E-016    $ (-2980 91.5 -2979.999 96.5)CMOSN560 88 88 D_lateral AREA=3.125E-016    
* Pins of element D559 are shorted:
* D559 104 104 D_lateral AREA=3.125E-016    $ (-2922.5 121.999 -2917.5 122)CMOSN559 104 104 D_lateral AREA=3.125E-016    
* Pins of element D558 are shorted:
* D558 104 104 D_lateral AREA=3.125E-016    $ (-2916 77.999 -2911 78)CMOSN558 104 104 D_lateral AREA=3.125E-016    
M557 2668 2470 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M556 88 2495 2470 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M555 2461 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M553 2464 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M552 2464 2463 2461 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M551 2462 2197 2457 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M550 2462 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D549 are shorted:
* D549 88 88 D_lateral AREA=3.125E-016    $ (-3080.5 91.5 -3080.499 96.5)CMOSN549 88 88 D_lateral AREA=3.125E-016    
M548 88 2666 2489 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M547 2666 2667 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M546 2470 2467 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M545 88 2467 2667 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M544 2667 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M543 2478 2480 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M542 2466 2074 2467 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M541 2467 2471 2472 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M540 2471 2485 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M539 104 2074 2465 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M538 2472 2465 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M537 104 2485 2466 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M536 104 2666 2486 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M535 2666 2667 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M534 104 2470 2668 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M533 2469 2467 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M532 2470 2495 2469 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M531 2667 2467 2468 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M530 2468 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M529 2478 2480 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D527 are shorted:
* D527 104 104 D_lateral AREA=3.125E-016    $ (-3163.5 121.999 -3158.5 122)CMOSN527 104 104 D_lateral AREA=3.125E-016    
* Pins of element D526 are shorted:
* D526 88 88 D_lateral AREA=3.125E-016    $ (-3174.5 46.5 -3174.499 51.5)CMOSN526 88 88 D_lateral AREA=3.125E-016    
* Pins of element D525 are shorted:
* D525 104 104 D_lateral AREA=3.125E-016    $ (-3173.001 29.5 -3173 34.5)CMOSN525 104 104 D_lateral AREA=3.125E-016    
* Pins of element D524 are shorted:
* D524 88 88 D_lateral AREA=3.125E-016    $ (-3125 91.5 -3124.999 96.5)CMOSN524 88 88 D_lateral AREA=3.125E-016    
M523 2525 2486 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M522 2489 2668 2490 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M521 2490 2492 2486 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M520 88 2478 2476 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M519 88 2478 2488 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M518 2488 2475 2498 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M517 2475 2479 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M516 2487 2479 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M515 2498 2476 2487 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M514 2525 2486 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M513 2486 2668 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M512 104 2492 2486 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M511 2474 2485 2479 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M510 2479 2483 2484 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M509 2483 2491 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M508 104 2485 2473 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M507 2484 2473 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M506 104 2491 2474 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M505 2482 2197 2480 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M504 2482 2495 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M503 2477 2478 2498 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M502 104 2478 2476 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M501 2498 2475 2481 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M500 104 2479 2477 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M499 2475 2479 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M498 2481 2476 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D496 are shorted:
* D496 88 88 D_lateral AREA=3.125E-016    $ (-3219 91.999 -3214 92)CMOSN496 88 88 D_lateral AREA=3.125E-016    
* Pins of element D495 are shorted:
* D495 104 104 D_lateral AREA=3.125E-016    $ (-3287.5 77.999 -3282.5 78)CMOSN495 104 104 D_lateral AREA=3.125E-016    
M494 2492 2493 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M493 88 2495 2493 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M492 2493 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M491 104 2494 2491 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M490 2492 2493 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M489 2493 2495 2497 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M488 2497 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M487 2494 2197 2496 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M486 2496 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D485 are shorted:
* D485 88 88 D_lateral AREA=3.125E-016    $ (-3351.5 91.5 -3351.499 96.5)CMOSN485 88 88 D_lateral AREA=3.125E-016    
* Pins of element D484 are shorted:
* D484 104 104 D_lateral AREA=3.125E-016    $ (-3294 121.999 -3289 122)CMOSN484 104 104 D_lateral AREA=3.125E-016    
M483 2670 2669 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M482 88 2525 2669 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M481 2669 2506 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M480 2500 2074 2506 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M479 104 2074 2505 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M478 2670 2669 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M477 2669 2525 2499 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M476 2499 2506 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D475 are shorted:
* D475 88 88 D_lateral AREA=3.125E-016    $ (-3453 91.5 -3452.999 96.5)CMOSN475 88 88 D_lateral AREA=3.125E-016    
M474 2508 2670 2509 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M473 88 2671 2508 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M472 2509 2516 2673 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M471 2671 2672 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M470 88 2506 2672 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M469 2672 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M468 2515 2502 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M467 2506 2501 2507 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M466 2501 2165 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M465 2507 2505 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M464 104 2165 2500 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M463 2673 2670 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M462 104 2671 2673 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M461 104 2516 2673 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M460 2671 2672 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M459 2672 2506 2504 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M458 2504 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M457 2515 2502 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M456 2502 2197 2503 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M455 2503 2525 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D453 are shorted:
* D453 104 104 D_lateral AREA=3.125E-016    $ (-3536 121.999 -3531 122)CMOSN453 104 104 D_lateral AREA=3.125E-016    
* Pins of element D452 are shorted:
* D452 104 104 D_lateral AREA=3.125E-016    $ (-3545.501 29.5 -3545.5 34.5)CMOSN452 104 104 D_lateral AREA=3.125E-016    
* Pins of element D451 are shorted:
* D451 88 88 D_lateral AREA=3.125E-016    $ (-3547 46.5 -3546.999 51.5)CMOSN451 88 88 D_lateral AREA=3.125E-016    
* Pins of element D450 are shorted:
* D450 88 88 D_lateral AREA=3.125E-016    $ (-3497.5 91.5 -3497.499 96.5)CMOSN450 88 88 D_lateral AREA=3.125E-016    
M448 2677 2673 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M447 2516 2524 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M446 88 2515 2513 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M445 88 2515 2523 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M444 2523 2512 2529 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M443 2512 2517 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M442 2522 2517 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M441 2529 2513 2522 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M440 2677 2673 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M439 2516 2524 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M438 2511 2165 2517 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M437 2517 2520 2521 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M436 2520 2519 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M435 104 2165 2510 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M434 2521 2510 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M433 104 2519 2511 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M432 2514 2515 2529 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M431 2513 2515 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M430 2529 2512 2518 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M429 104 2517 2514 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M428 2512 2517 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M427 2518 2513 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D426 are shorted:
* D426 104 104 D_lateral AREA=3.125E-016    $ (-3666.5 121.999 -3661.5 122)CMOSN426 104 104 D_lateral AREA=3.125E-016    
* Pins of element D425 are shorted:
* D425 88 88 D_lateral AREA=3.125E-016    $ (-3591.5 91.999 -3586.5 92)CMOSN425 88 88 D_lateral AREA=3.125E-016    
* Pins of element D424 are shorted:
* D424 104 104 D_lateral AREA=3.125E-016    $ (-3660 77.999 -3655 78)CMOSN424 104 104 D_lateral AREA=3.125E-016    
M423 88 2525 2524 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M422 2524 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M421 104 2526 2519 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M420 2524 2525 2528 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M419 2528 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M418 2526 2197 2527 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M417 2527 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D416 are shorted:
* D416 88 88 D_lateral AREA=3.125E-016    $ (-3724 91.5 -3723.999 96.5)CMOSN416 88 88 D_lateral AREA=3.125E-016    
M415 88 2074 2675 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M414 88 2074 2537 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M413 2537 2674 2545 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M412 2674 2678 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M411 2536 2678 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M410 2545 2675 2536 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M409 2074 2531 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M408 88 2180 2531 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M407 2531 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M406 2530 2074 2545 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M405 2675 2074 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M404 2545 2674 2535 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M403 2530 2678 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M402 2674 2678 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M401 2535 2675 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M400 2074 2531 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M399 2531 2180 2534 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M398 2534 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M397 2197 2533 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M396 104 2532 2533 104 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M395 2533 491 104 104 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
* Pins of element D394 are shorted:
* D394 88 88 D_lateral AREA=3.125E-016    $ (-3921 45.499 -3916 45.5)CMOSN394 88 88 D_lateral AREA=3.125E-016    
* Pins of element D393 are shorted:
* D393 104 104 D_lateral AREA=3.125E-016    $ (-3989.5 31.499 -3984.5 31.5)CMOSN393 104 104 D_lateral AREA=3.125E-016    
* Pins of element D392 are shorted:
* D392 88 88 D_lateral AREA=3.125E-016    $ (-3944 90 -3943.999 95)CMOSN392 88 88 D_lateral AREA=3.125E-016    
M391 2678 2676 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M390 88 2677 2676 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M389 2676 491 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M388 2532 2538 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M387 88 2540 2538 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M386 2538 2539 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M385 2539 491 88 88 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M384 2678 2676 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M383 2676 2677 2544 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M382 2544 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M381 2532 2538 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M380 2538 2540 2543 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M379 2543 2539 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M378 2539 491 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M377 2201 2542 104 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M376 2542 2540 2541 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M375 2541 491 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D374 are shorted:
* D374 88 88 D_lateral AREA=3.125E-016    $ (-4049 45 -4048.999 50)CMOSN374 88 88 D_lateral AREA=3.125E-016    
* Pins of element D373 are shorted:
* D373 88 88 D_lateral AREA=3.125E-016    $ (-4028 90 -4027.999 95)CMOSN373 88 88 D_lateral AREA=3.125E-016    
* Pins of element D371 are shorted:
* D371 88 88 D_lateral AREA=3.125E-016    $ (216.5 -71 216.501 -66)CMOSN371 88 88 D_lateral AREA=3.125E-016    
M370 88 104 2547 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M369 88 104 2554 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M368 2554 2546 2682 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M367 2546 2211 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M366 2553 2211 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M365 2682 2547 2553 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M364 2681 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M363 2681 2682 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M362 88 2682 2680 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M361 2680 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M360 2688 2691 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M358 2548 104 2682 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M357 104 104 2547 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M356 2682 2546 2552 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M355 104 2211 2548 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M354 2546 2211 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M353 2552 2547 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D352 are shorted:
* D352 88 88 D_lateral AREA=3.125E-016    $ (202 -26.501 207 -26.5)CMOSN352 88 88 D_lateral AREA=3.125E-016    
* Pins of element D351 are shorted:
* D351 104 104 D_lateral AREA=3.125E-016    $ (133.5 -40.501 138.5 -40.5)CMOSN351 104 104 D_lateral AREA=3.125E-016    
* Pins of element D350 are shorted:
* D350 88 88 D_lateral AREA=3.125E-016    $ (172 -71 172.001 -66)CMOSN350 88 88 D_lateral AREA=3.125E-016    
* Pins of element D349 are shorted:
* D349 88 88 D_lateral AREA=3.125E-016    $ (117.5 -27 117.501 -22)CMOSN349 88 88 D_lateral AREA=3.125E-016    
M348 88 2211 2556 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M347 88 2211 2566 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M346 2566 2555 2697 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M345 2555 2568 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M344 2565 2568 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M343 2697 2556 2565 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M342 2691 2564 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M341 2691 104 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M340 88 2688 2686 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M339 88 2688 2563 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M338 2685 2697 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M337 2563 2685 2699 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M336 2562 2697 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M335 2699 2686 2562 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M334 2557 2211 2697 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M333 104 2211 2556 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M332 2697 2555 2561 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M331 104 2568 2557 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M330 2555 2568 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M329 2561 2556 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M328 2691 2564 2560 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M327 2560 104 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D326 are shorted:
* D326 88 88 D_lateral AREA=3.125E-016    $ (71.5 -26.501 76.5 -26.5)CMOSN326 88 88 D_lateral AREA=3.125E-016    
* Pins of element D325 are shorted:
* D325 88 88 D_lateral AREA=3.125E-016    $ (78 -70.501 83 -70.5)CMOSN325 88 88 D_lateral AREA=3.125E-016    
M324 88 2567 2568 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M323 2695 2696 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M322 88 104 2696 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M321 2696 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M320 88 2564 2567 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M319 2567 103 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M318 104 2567 2568 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M317 2567 2564 2569 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M316 2569 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D315 are shorted:
* D315 88 88 D_lateral AREA=3.125E-016    $ (-54.5 -71 -54.499 -66)CMOSN315 88 88 D_lateral AREA=3.125E-016    
* Pins of element D314 are shorted:
* D314 104 104 D_lateral AREA=3.125E-016    $ (3 -40.501 8 -40.5)CMOSN314 104 104 D_lateral AREA=3.125E-016    
* Pins of element D313 are shorted:
* D313 88 88 D_lateral AREA=3.125E-016    $ (-54 -27 -53.999 -22)CMOSN313 88 88 D_lateral AREA=3.125E-016    
M312 88 104 2580 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M311 88 104 2571 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M310 2571 2577 2579 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M309 88 2717 2700 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M308 2700 2579 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M307 2572 104 2579 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M306 104 104 2580 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D305 are shorted:
* D305 88 88 D_lateral AREA=3.125E-016    $ (-161.5 -26.501 -156.5 -26.5)CMOSN305 88 88 D_lateral AREA=3.125E-016    
* Pins of element D304 are shorted:
* D304 88 88 D_lateral AREA=3.125E-016    $ (-147 -71 -146.999 -66)CMOSN304 88 88 D_lateral AREA=3.125E-016    
M303 2577 2238 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M302 2581 2238 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M301 2579 2580 2581 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M300 88 2579 2704 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M299 2704 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M298 2587 2705 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M297 88 2564 2705 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M296 2705 2717 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M295 2710 2587 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M294 2579 2577 2578 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M293 104 2238 2572 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M292 2577 2238 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M291 2578 2580 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M289 2705 2564 2576 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M288 2576 2717 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D287 are shorted:
* D287 104 104 D_lateral AREA=3.125E-016    $ (-230 -40.501 -225 -40.5)CMOSN287 104 104 D_lateral AREA=3.125E-016    
* Pins of element D286 are shorted:
* D286 88 88 D_lateral AREA=3.125E-016    $ (-191.5 -71 -191.499 -66)CMOSN286 88 88 D_lateral AREA=3.125E-016    
* Pins of element D284 are shorted:
* D284 88 88 D_lateral AREA=3.125E-016    $ (-246 -27 -245.999 -22)CMOSN284 88 88 D_lateral AREA=3.125E-016    
* Pins of element D283 are shorted:
* D283 88 88 D_lateral AREA=3.125E-016    $ (-285.5 -70.501 -280.5 -70.5)CMOSN283 88 88 D_lateral AREA=3.125E-016    
M282 88 2591 2592 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M281 2713 2716 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M280 88 2238 2583 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M279 88 2238 2590 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M278 2590 2582 2714 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M277 2582 2592 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M276 2589 2592 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M275 2714 2583 2589 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M274 88 2587 2588 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M273 2711 2714 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M272 2588 2711 2722 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M271 2586 2714 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M270 2722 2710 2586 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M269 104 2591 2592 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M268 2584 2238 2714 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M267 2583 2238 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M266 2714 2582 2585 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M265 104 2592 2584 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M264 2582 2592 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M263 2585 2583 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D262 are shorted:
* D262 88 88 D_lateral AREA=3.125E-016    $ (-292 -26.501 -287 -26.5)CMOSN262 88 88 D_lateral AREA=3.125E-016    
* Pins of element D261 are shorted:
* D261 104 104 D_lateral AREA=3.125E-016    $ (-360.5 -40.501 -355.5 -40.5)CMOSN261 104 104 D_lateral AREA=3.125E-016    
M260 88 2717 2716 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M259 2716 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M258 88 2564 2591 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M257 2591 123 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M256 2591 2564 2593 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M255 2593 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D254 are shorted:
* D254 88 88 D_lateral AREA=3.125E-016    $ (-418 -71 -417.999 -66)CMOSN254 88 88 D_lateral AREA=3.125E-016    
* Pins of element D253 are shorted:
* D253 88 88 D_lateral AREA=3.125E-016    $ (-417.5 -27 -417.499 -22)CMOSN253 88 88 D_lateral AREA=3.125E-016    
M252 88 104 2595 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M251 88 104 2601 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M250 2601 2594 2721 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M249 2594 2270 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M248 2600 2270 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M247 2721 2595 2600 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M246 88 2740 2720 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M245 2720 2721 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M244 88 2721 2719 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M243 2719 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M242 2596 104 2721 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M241 104 104 2595 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M240 2721 2594 2599 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M239 104 2270 2596 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M238 2594 2270 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M237 2599 2595 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D236 are shorted:
* D236 88 88 D_lateral AREA=3.125E-016    $ (-526 -26.501 -521 -26.5)CMOSN236 88 88 D_lateral AREA=3.125E-016    
* Pins of element D234 are shorted:
* D234 88 88 D_lateral AREA=3.125E-016    $ (-511.5 -71 -511.499 -66)CMOSN234 88 88 D_lateral AREA=3.125E-016    
* Pins of element D233 are shorted:
* D233 88 88 D_lateral AREA=3.125E-016    $ (-556 -71 -555.999 -66)CMOSN233 88 88 D_lateral AREA=3.125E-016    
M232 2726 2729 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M231 88 2270 2613 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M230 88 2270 2608 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M229 2608 2609 2612 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M228 88 2564 2729 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M227 2729 2740 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M226 88 2726 2725 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M225 88 2726 2607 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M224 2607 2733 2737 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M222 2737 2725 2606 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M221 2610 2270 2612 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M220 104 2270 2613 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M219 2612 2609 2605 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M217 2729 2564 2604 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M216 2604 2740 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D215 are shorted:
* D215 104 104 D_lateral AREA=3.125E-016    $ (-594.5 -40.501 -589.5 -40.5)CMOSN215 104 104 D_lateral AREA=3.125E-016    
* Pins of element D214 are shorted:
* D214 88 88 D_lateral AREA=3.125E-016    $ (-656.5 -26.501 -651.5 -26.5)CMOSN214 88 88 D_lateral AREA=3.125E-016    
* Pins of element D213 are shorted:
* D213 88 88 D_lateral AREA=3.125E-016    $ (-610.5 -27 -610.499 -22)CMOSN213 88 88 D_lateral AREA=3.125E-016    
* Pins of element D212 are shorted:
* D212 88 88 D_lateral AREA=3.125E-016    $ (-650 -70.501 -645 -70.5)CMOSN212 88 88 D_lateral AREA=3.125E-016    
M211 88 2615 2611 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M210 2735 2738 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M208 2609 2611 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M207 2614 2611 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M206 2612 2613 2614 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M205 88 2564 2615 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M204 2733 2612 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M203 88 2612 2606 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M202 104 2615 2611 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M201 2609 2611 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M200 104 2611 2610 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M199 104 2613 2605 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=187.5f PS=1.25u    
* Pins of element D198 are shorted:
* D198 88 88 D_lateral AREA=3.125E-016    $ (-782.5 -71 -782.499 -66)CMOSN198 88 88 D_lateral AREA=3.125E-016    
* Pins of element D197 are shorted:
* D197 104 104 D_lateral AREA=3.125E-016    $ (-725 -40.501 -720 -40.5)CMOSN197 104 104 D_lateral AREA=3.125E-016    
* Pins of element D196 are shorted:
* D196 88 88 D_lateral AREA=3.125E-016    $ (-782 -27 -781.999 -22)CMOSN196 88 88 D_lateral AREA=3.125E-016    
M195 2738 2740 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M194 2738 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M193 2615 145 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M191 88 2760 2744 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M189 2615 2564 2616 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M188 2616 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M187 104 104 2618 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D186 are shorted:
* D186 88 88 D_lateral AREA=3.125E-016    $ (-889.5 -26.501 -884.5 -26.5)CMOSN186 88 88 D_lateral AREA=3.125E-016    
* Pins of element D185 are shorted:
* D185 88 88 D_lateral AREA=3.125E-016    $ (-875 -71 -874.999 -66)CMOSN185 88 88 D_lateral AREA=3.125E-016    
M184 2618 104 88 88 CMOSP L=500n W=750n AD=2p PD=6u AS=1.90625p PS=5.75u    
M183 88 104 2626 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M182 2626 2617 2745 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M181 2617 2308 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M180 2625 2308 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M179 2745 2618 2625 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M178 88 2745 2744 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M177 88 2745 2743 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M176 2743 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M175 2752 2746 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M174 88 2564 2746 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M172 2619 104 2745 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M171 2745 2617 2624 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M170 104 2308 2619 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M169 2617 2308 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M168 2624 2618 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M167 2746 2564 2623 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
* Pins of element D165 are shorted:
* D165 104 104 D_lateral AREA=3.125E-016    $ (-958 -40.501 -953 -40.5)CMOSN165 104 104 D_lateral AREA=3.125E-016    
* Pins of element D164 are shorted:
* D164 88 88 D_lateral AREA=3.125E-016    $ (-919.5 -71 -919.499 -66)CMOSN164 88 88 D_lateral AREA=3.125E-016    
* Pins of element D163 are shorted:
* D163 88 88 D_lateral AREA=3.125E-016    $ (-974 -27 -973.999 -22)CMOSN163 88 88 D_lateral AREA=3.125E-016    
M162 88 2308 2628 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M161 88 2308 2635 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M160 2635 2627 2755 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M159 2627 2637 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M158 2634 2637 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M157 2755 2628 2634 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M156 88 2760 2746 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M155 88 2752 2750 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=2p PS=6u    
M154 88 2752 2633 88 CMOSP L=500n W=750n AD=1.90625p PD=5.75u AS=187.5f PS=1.25u    
M153 2749 2755 88 88 CMOSP L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M152 2633 2749 2762 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.9453125p PS=4.5u    
M151 2632 2755 88 88 CMOSP L=500n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M150 2762 2750 2632 88 CMOSP L=500n W=750n AD=1.9453125p PD=4.5u AS=187.5f PS=1.25u    
M149 2629 2308 2755 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M148 104 2308 2628 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M147 2755 2627 2631 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M146 104 2637 2629 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M145 2627 2637 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M144 2631 2628 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
M143 104 2760 2623 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
* Pins of element D142 are shorted:
* D142 88 88 D_lateral AREA=3.125E-016    $ (-1020 -26.501 -1015 -26.5)CMOSN142 88 88 D_lateral AREA=3.125E-016    
* Pins of element D141 are shorted:
* D141 104 104 D_lateral AREA=3.125E-016    $ (-1088.5 -40.501 -1083.5 -40.5)CMOSN141 104 104 D_lateral AREA=3.125E-016    
* Pins of element D140 are shorted:
* D140 88 88 D_lateral AREA=3.125E-016    $ (-1013.5 -70.501 -1008.5 -70.5)CMOSN140 88 88 D_lateral AREA=3.125E-016    
M139 88 2636 2637 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M138 2758 2759 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M137 88 2760 2759 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M136 2759 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M135 88 2564 2636 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M134 2636 167 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M133 104 2636 2637 104 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M132 2636 2564 2638 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M131 2638 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D130 are shorted:
* D130 88 88 D_lateral AREA=3.125E-016    $ (-1146 -71 -1145.999 -66)CMOSN130 88 88 D_lateral AREA=3.125E-016    
* Pins of element D129 are shorted:
* D129 88 88 D_lateral AREA=3.125E-016    $ (-1145.5 -27 -1145.499 -22)CMOSN129 88 88 D_lateral AREA=3.125E-016    
M128 88 491 2641 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M127 2564 2641 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M126 2564 2641 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D125 are shorted:
* D125 88 88 D_lateral AREA=3.125E-016    $ (-1281.5 -27 -1281.499 -22)CMOSN125 88 88 D_lateral AREA=3.125E-016    
M124 2642 2545 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M123 2641 2642 88 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M122 2642 2545 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M121 2644 2642 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M120 2641 491 2644 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M119 88 2679 2693 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M118 2679 2680 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M117 2690 2681 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M116 104 2679 2689 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M115 2679 2680 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M114 2690 2681 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M113 2681 104 2684 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M112 2684 2682 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M111 2680 2682 2683 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M110 2683 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M109 2688 2691 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D108 are shorted:
* D108 88 88 D_lateral AREA=3.125E-016    $ (122.5 -116 122.501 -111)CMOSN108 88 88 D_lateral AREA=3.125E-016    
* Pins of element D107 are shorted:
* D107 104 104 D_lateral AREA=3.125E-016    $ (123.999 -133 124 -128)CMOSN107 104 104 D_lateral AREA=3.125E-016    
M106 2717 2689 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M105 2693 2690 2694 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M104 2694 2695 2689 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M103 2717 2689 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M102 2689 2690 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M101 104 2695 2689 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M100 2687 2688 2699 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M99 104 2688 2686 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M98 2699 2685 2692 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M97 104 2697 2687 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M96 2685 2697 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M95 2692 2686 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D94 are shorted:
* D94 104 104 D_lateral AREA=3.125E-016    $ (9.5 -84.501 14.5 -84.5)CMOSN94 104 104 D_lateral AREA=3.125E-016    
M93 2695 2696 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M92 2696 104 2698 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M91 2698 103 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M90 2702 2700 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M89 2702 2700 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M88 2700 2717 2701 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M87 2701 2579 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M86 2707 2702 2708 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M85 88 2703 2707 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M84 2708 2713 2709 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M83 2703 2704 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M82 2709 2702 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M81 104 2703 2709 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M80 104 2713 2709 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M79 2703 2704 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M78 2704 2579 2706 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M77 2706 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M76 2587 2705 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M75 104 2587 2710 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
* Pins of element D74 are shorted:
* D74 104 104 D_lateral AREA=3.125E-016    $ (-239.501 -133 -239.5 -128)CMOSN74 104 104 D_lateral AREA=3.125E-016    
* Pins of element D73 are shorted:
* D73 88 88 D_lateral AREA=3.125E-016    $ (-241 -116 -240.999 -111)CMOSN73 88 88 D_lateral AREA=3.125E-016    
M72 2740 2709 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M71 2740 2709 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M70 2713 2716 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M69 2712 2587 2722 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M68 2722 2711 2715 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M67 104 2714 2712 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M66 2711 2714 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M65 2715 2710 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D64 are shorted:
* D64 104 104 D_lateral AREA=3.125E-016    $ (-354 -84.501 -349 -84.5)CMOSN64 104 104 D_lateral AREA=3.125E-016    
M63 2716 2717 2718 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M62 2718 123 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M61 2728 2719 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M60 2727 2720 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M59 2728 2719 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M58 2727 2720 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M57 2720 2740 2724 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M56 2724 2721 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M55 2719 2721 2723 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M54 2723 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M53 2760 2736 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M52 2731 2727 2732 88 CMOSP L=750n W=750n AD=1.125p PD=3.75u AS=796.875f PS=2.875u    
M51 88 2728 2731 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M50 2732 2735 2736 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M49 2760 2736 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M48 2736 2727 104 104 CMOSN L=1.5u W=750n AD=1.15625p PD=3.5u AS=1.203125p PS=3.375u    
M47 104 2728 2736 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M46 104 2735 2736 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M45 2726 2729 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M44 2734 2726 2737 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M43 104 2726 2725 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M42 2737 2733 2730 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M41 2730 2725 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D40 are shorted:
* D40 104 104 D_lateral AREA=3.125E-016    $ (-604.001 -133 -604 -128)CMOSN40 104 104 D_lateral AREA=3.125E-016    
* Pins of element D39 are shorted:
* D39 88 88 D_lateral AREA=3.125E-016    $ (-605.5 -116 -605.499 -111)CMOSN39 88 88 D_lateral AREA=3.125E-016    
M38 2735 2738 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M37 2733 2612 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M36 104 2612 2734 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D35 are shorted:
* D35 104 104 D_lateral AREA=3.125E-016    $ (-718.5 -84.501 -713.5 -84.5)CMOSN35 104 104 D_lateral AREA=3.125E-016    
M34 2754 2744 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M33 2738 2740 2741 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M32 2741 145 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M31 2754 2744 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M30 2744 2760 2739 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M27 88 2742 2748 88 CMOSP L=750n W=750n AD=1.59375p PD=5.25u AS=1.125p PS=3.75u    
M26 2742 2743 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M24 104 2742 2753 104 CMOSN L=1.5u W=750n AD=1.59375p PD=5.25u AS=1.15625p PS=3.5u    
M23 2742 2743 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M22 104 2745 2739 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M21 2743 2745 2747 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M20 2747 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M19 2752 2746 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
* Pins of element D18 are shorted:
* D18 88 88 D_lateral AREA=3.125E-016    $ (-969 -116 -968.999 -111)CMOSN18 88 88 D_lateral AREA=3.125E-016    
* Pins of element D17 are shorted:
* D17 104 104 D_lateral AREA=3.125E-016    $ (-967.501 -133 -967.5 -128)CMOSN17 104 104 D_lateral AREA=3.125E-016    
M16 2763 2753 88 88 CMOSP L=500n W=2u AD=3.0625p PD=8u AS=3.0625p PS=8u    
M15 2757 2754 2748 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.125p PS=3.75u    
M14 2757 2758 2753 88 CMOSP L=750n W=750n AD=796.875f PD=2.875u AS=1.75p PS=5.5u    
M13 2763 2753 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M12 104 2754 2753 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=1.15625p PS=3.5u    
M11 104 2758 2753 104 CMOSN L=1.5u W=750n AD=1.203125p PD=3.375u AS=3.15625p PS=9.25u    
M10 2751 2752 2762 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.84375p PS=4.375u    
M9 104 2752 2750 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M8 2762 2749 2756 104 CMOSN L=500n W=750n AD=1.84375p PD=4.375u AS=187.5f PS=1.25u    
M7 104 2755 2751 104 CMOSN L=500n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M6 2749 2755 104 104 CMOSN L=500n W=750n AD=1.75p PD=5.5u AS=2.21875p PS=6.25u    
M5 2756 2750 104 104 CMOSN L=500n W=750n AD=187.5f PD=1.25u AS=968.75f PS=3u    
* Pins of element D4 are shorted:
* D4 104 104 D_lateral AREA=3.125E-016    $ (-1082 -84.501 -1077 -84.5)CMOSN4 104 104 D_lateral AREA=3.125E-016    
M3 2758 2759 104 104 CMOSN L=750n W=750n AD=2.03125p PD=6.25u AS=2.03125p PS=6.25u    
M2 2759 2760 2761 104 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1 2761 167 104 104 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    

* Total Nodes: 2763
* Total Elements: 5977
* Total Number of Shorted Elements not written to the SPICE file: 0
* Output Generation Elapsed Time: 7.078 sec
* Total Extract Elapsed Time: 22.250 sec

* INPUTS 
VVDD 88 0 5v
VGND 104 0 0v
VLf7 183 0 0v
VLf6 357 0 0v
VLf5 664 0 0v
VLf4 973 0 0v
VLf3 1269 0 0v
VLf2 1484 0 0v
VLf1 2177 0 0v
VLf0 2540 0 0v
VZ 491 0 5v
VBf3 167 0 5v
VBf2 145 0 5v
VBf1 123 0 5v
VBf0 103 0 5v

* OUTPUTS 
*Q0 2545
*Q1 2180
*Q2 2017
*Q3 1481
*Q4 976
*Q5 819
*Q6 482
*Q7 186
*r0 2699
*r1 2722
*r2 2737
*r3 2762
*Sf4 2335
*Sf5 2368
*Sf6 2403
*Sf7 2428
* OUTPUT can be put in trace in simulation 
*  V(2545) V(2180) V(2017) V(1481) V(976) V(819) V(482) V(186) V(2699) V(2722) V(2737) V(2762) V(2335) V(2368) V(2403) V(2428)
.op
.tran 0.1ns 100ns
.probe
.END